// ============================================================================
// Amazon FPGA Hardware Development Kit
//
// Copyright 2024 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
// ============================================================================


//====================================================================================
// Top level module file for prospero
//====================================================================================

module prospero
    #(
      parameter EN_DDR = 0,
      parameter EN_HBM = 0
    )
    (
      `include "cl_ports.vh"
    );

`include "cl_id_defines.vh" // CL ID defines required for all examples
`include "prospero_defines.vh"


//=============================================================================
// GLOBALS
//=============================================================================

  always_comb begin
     cl_sh_flr_done    = 'b1;
     cl_sh_status0     = 'b0;
     cl_sh_status1     = 'b0;
     cl_sh_status2     = 'b0;
     cl_sh_id0         = `CL_SH_ID0;
     cl_sh_id1         = `CL_SH_ID1;
     cl_sh_status_vled = 'b0;
     cl_sh_dma_wr_full = 'b0;
     cl_sh_dma_rd_full = 'b0;
  end

//=============================================================================
// Circuit Instance and Registers
//=============================================================================

  // Parameters for the circuit
  localparam CIRCUIT_WIDTH = 64;
  localparam CIRCUIT_FRAC_BITS = 32;
  
  // Registers to store inputs and outputs
  logic [CIRCUIT_WIDTH-1:0] reg_x;
  logic [CIRCUIT_WIDTH-1:0] reg_y;
  logic [CIRCUIT_WIDTH-1:0] reg_out;
  
  // Circuit instance
  circuit_wrapper #(
    .WIDTH(CIRCUIT_WIDTH),
    .FRAC_BITS(CIRCUIT_FRAC_BITS)
  ) circuit_wrapper_inst (
    .clk(clk_main_a0),
    .reset(~rst_main_n),
    .x(reg_x_pipe),
    .y(reg_y_pipe),
    .out(reg_out_pipe)
  );

//=============================================================================
// PCIM
//=============================================================================

  // Cause Protocol Violations
  always_comb begin
    cl_sh_pcim_awaddr  = 'b0;
    cl_sh_pcim_awsize  = 'b0;
    cl_sh_pcim_awburst = 'b0;
    cl_sh_pcim_awvalid = 'b0;

    cl_sh_pcim_wdata   = 'b0;
    cl_sh_pcim_wstrb   = 'b0;
    cl_sh_pcim_wlast   = 'b0;
    cl_sh_pcim_wvalid  = 'b0;

    cl_sh_pcim_araddr  = 'b0;
    cl_sh_pcim_arsize  = 'b0;
    cl_sh_pcim_arburst = 'b0;
    cl_sh_pcim_arvalid = 'b0;
  end

  // Remaining CL Output Ports
  always_comb begin
    cl_sh_pcim_awid    = 'b0;
    cl_sh_pcim_awlen   = 'b0;
    cl_sh_pcim_awcache = 'b0;
    cl_sh_pcim_awlock  = 'b0;
    cl_sh_pcim_awprot  = 'b0;
    cl_sh_pcim_awqos   = 'b0;
    cl_sh_pcim_awuser  = 'b0;

    cl_sh_pcim_wid     = 'b0;
    cl_sh_pcim_wuser   = 'b0;

    cl_sh_pcim_arid    = 'b0;
    cl_sh_pcim_arlen   = 'b0;
    cl_sh_pcim_arcache = 'b0;
    cl_sh_pcim_arlock  = 'b0;
    cl_sh_pcim_arprot  = 'b0;
    cl_sh_pcim_arqos   = 'b0;
    cl_sh_pcim_aruser  = 'b0;

    cl_sh_pcim_rready  = 'b0;
  end

//=============================================================================
// PCIS
//=============================================================================

  // Cause Protocol Violations
  always_comb begin
    cl_sh_dma_pcis_bresp   = 'b0;
    cl_sh_dma_pcis_rresp   = 'b0;
    cl_sh_dma_pcis_rvalid  = 'b0;
  end

  // Remaining CL Output Ports
  always_comb begin
    cl_sh_dma_pcis_awready = 'b0;

    cl_sh_dma_pcis_wready  = 'b0;

    cl_sh_dma_pcis_bid     = 'b0;
    cl_sh_dma_pcis_bvalid  = 'b0;

    cl_sh_dma_pcis_arready  = 'b0;

    cl_sh_dma_pcis_rid     = 'b0;
    cl_sh_dma_pcis_rdata   = 'b0;
    cl_sh_dma_pcis_rlast   = 'b0;
    cl_sh_dma_pcis_ruser   = 'b0;
  end

//=============================================================================
// OCL - Interface for CPU Communication with Circuit
//=============================================================================

  // Address decoding for register access via OCL AXI-Lite
  localparam REG_X_ADDR_LOW     = 32'h00;  // Address for x input (lower 32 bits)
  localparam REG_X_ADDR_HIGH    = 32'h04;  // Address for x input (upper 32 bits)
  localparam REG_Y_ADDR_LOW     = 32'h08;  // Address for y input (lower 32 bits)
  localparam REG_Y_ADDR_HIGH    = 32'h0C;  // Address for y input (upper 32 bits)
  localparam REG_OUT_ADDR_LOW   = 32'h10;  // Address for circuit output (lower 32 bits)
  localparam REG_OUT_ADDR_HIGH  = 32'h14;  // Address for circuit output (upper 32 bits)

  // Registers for OCL AXI-Lite response
  logic [31:0] ocl_read_data;
  logic ocl_read_valid;
  logic ocl_write_valid;
  
  // AXI-Lite write logic
  always_ff @(posedge clk_main_a0) begin
    if (!rst_main_n) begin
      reg_x <= 0;
      reg_y <= 0;
      ocl_write_valid <= 1'b0;
    end else begin
      ocl_write_valid <= 1'b0;
      
      if (ocl_cl_awvalid && ocl_cl_wvalid) begin
        ocl_write_valid <= 1'b1;
        
        case (ocl_cl_awaddr[7:0])
          REG_X_ADDR_LOW:  reg_x[31:0]  <= ocl_cl_wdata;
          REG_X_ADDR_HIGH: reg_x[63:32] <= ocl_cl_wdata;
          REG_Y_ADDR_LOW:  reg_y[31:0]  <= ocl_cl_wdata;
          REG_Y_ADDR_HIGH: reg_y[63:32] <= ocl_cl_wdata;
          default: ; // No operation
        endcase
      end
    end
  end
  
  // AXI-Lite read logic
  always_ff @(posedge clk_main_a0) begin
    if (!rst_main_n) begin
      ocl_read_data <= 0;
      ocl_read_valid <= 1'b0;
    end else begin
      ocl_read_valid <= 1'b0;
      
      if (ocl_cl_arvalid) begin
        ocl_read_valid <= 1'b1;
        
        case (ocl_cl_araddr[7:0])
          REG_X_ADDR_LOW:     ocl_read_data <= reg_x[31:0];
          REG_X_ADDR_HIGH:    ocl_read_data <= reg_x[63:32];
          REG_Y_ADDR_LOW:     ocl_read_data <= reg_y[31:0];
          REG_Y_ADDR_HIGH:    ocl_read_data <= reg_y[63:32];
          REG_OUT_ADDR_LOW:   ocl_read_data <= reg_out[31:0];
          REG_OUT_ADDR_HIGH:  ocl_read_data <= reg_out[63:32];
          default:            ocl_read_data <= 32'hDEADBEEF;
        endcase
      end
    end
  end

  // OCL AXI-Lite interface signals
  assign cl_ocl_awready = 1'b1;  // Always ready to accept write address
  assign cl_ocl_wready  = 1'b1;  // Always ready to accept write data
  assign cl_ocl_bvalid  = ocl_write_valid;
  assign cl_ocl_bresp   = 2'b00; // OKAY response
  
  assign cl_ocl_arready = 1'b1;  // Always ready to accept read address
  assign cl_ocl_rvalid  = ocl_read_valid;
  assign cl_ocl_rdata   = ocl_read_data;
  assign cl_ocl_rresp   = 2'b00; // OKAY response

//=============================================================================
// SDA
//=============================================================================

  // Cause Protocol Violations
  always_comb begin
    cl_sda_bresp   = 'b0;
    cl_sda_rresp   = 'b0;
    cl_sda_rvalid  = 'b0;
  end

  // Remaining CL Output Ports
  always_comb begin
    cl_sda_awready = 'b0;
    cl_sda_wready  = 'b0;

    cl_sda_bvalid = 'b0;

    cl_sda_arready = 'b0;

    cl_sda_rdata   = 'b0;
  end

//=============================================================================
// SH_DDR
//=============================================================================

   sh_ddr
     #(
       .DDR_PRESENT (EN_DDR)
       )
   SH_DDR
     (
      .clk                       (clk_main_a0 ),
      .rst_n                     (            ),
      .stat_clk                  (clk_main_a0 ),
      .stat_rst_n                (            ),
      .CLK_DIMM_DP               (CLK_DIMM_DP ),
      .CLK_DIMM_DN               (CLK_DIMM_DN ),
      .M_ACT_N                   (M_ACT_N     ),
      .M_MA                      (M_MA        ),
      .M_BA                      (M_BA        ),
      .M_BG                      (M_BG        ),
      .M_CKE                     (M_CKE       ),
      .M_ODT                     (M_ODT       ),
      .M_CS_N                    (M_CS_N      ),
      .M_CLK_DN                  (M_CLK_DN    ),
      .M_CLK_DP                  (M_CLK_DP    ),
      .M_PAR                     (M_PAR       ),
      .M_DQ                      (M_DQ        ),
      .M_ECC                     (M_ECC       ),
      .M_DQS_DP                  (M_DQS_DP    ),
      .M_DQS_DN                  (M_DQS_DN    ),
      .cl_RST_DIMM_N             (RST_DIMM_N  ),
      .cl_sh_ddr_axi_awid        (            ),
      .cl_sh_ddr_axi_awaddr      (            ),
      .cl_sh_ddr_axi_awlen       (            ),
      .cl_sh_ddr_axi_awsize      (            ),
      .cl_sh_ddr_axi_awvalid     (            ),
      .cl_sh_ddr_axi_awburst     (            ),
      .cl_sh_ddr_axi_awuser      (            ),
      .cl_sh_ddr_axi_awready     (            ),
      .cl_sh_ddr_axi_wdata       (            ),
      .cl_sh_ddr_axi_wstrb       (            ),
      .cl_sh_ddr_axi_wlast       (            ),
      .cl_sh_ddr_axi_wvalid      (            ),
      .cl_sh_ddr_axi_wready      (            ),
      .cl_sh_ddr_axi_bid         (            ),
      .cl_sh_ddr_axi_bresp       (            ),
      .cl_sh_ddr_axi_bvalid      (            ),
      .cl_sh_ddr_axi_bready      (            ),
      .cl_sh_ddr_axi_arid        (            ),
      .cl_sh_ddr_axi_araddr      (            ),
      .cl_sh_ddr_axi_arlen       (            ),
      .cl_sh_ddr_axi_arsize      (            ),
      .cl_sh_ddr_axi_arvalid     (            ),
      .cl_sh_ddr_axi_arburst     (            ),
      .cl_sh_ddr_axi_aruser      (            ),
      .cl_sh_ddr_axi_arready     (            ),
      .cl_sh_ddr_axi_rid         (            ),
      .cl_sh_ddr_axi_rdata       (            ),
      .cl_sh_ddr_axi_rresp       (            ),
      .cl_sh_ddr_axi_rlast       (            ),
      .cl_sh_ddr_axi_rvalid      (            ),
      .cl_sh_ddr_axi_rready      (            ),
      .sh_ddr_stat_bus_addr      (            ),
      .sh_ddr_stat_bus_wdata     (            ),
      .sh_ddr_stat_bus_wr        (            ),
      .sh_ddr_stat_bus_rd        (            ),
      .sh_ddr_stat_bus_ack       (            ),
      .sh_ddr_stat_bus_rdata     (            ),
      .ddr_sh_stat_int           (            ),
      .sh_cl_ddr_is_ready        (            )
      );

  always_comb begin
    cl_sh_ddr_stat_ack   = 'b0;
    cl_sh_ddr_stat_rdata = 'b0;
    cl_sh_ddr_stat_int   = 'b0;
  end

//=============================================================================
// USER-DEFIEND INTERRUPTS
//=============================================================================

  always_comb begin
    cl_sh_apppf_irq_req = 'b0;
  end

//=============================================================================
// VIRTUAL JTAG
//=============================================================================

  always_comb begin
    tdo = 'b0;
  end

//=============================================================================
// HBM MONITOR IO
//=============================================================================

  always_comb begin
    hbm_apb_paddr_1   = 'b0;
    hbm_apb_pprot_1   = 'b0;
    hbm_apb_psel_1    = 'b0;
    hbm_apb_penable_1 = 'b0;
    hbm_apb_pwrite_1  = 'b0;
    hbm_apb_pwdata_1  = 'b0;
    hbm_apb_pstrb_1   = 'b0;
    hbm_apb_pready_1  = 'b0;
    hbm_apb_prdata_1  = 'b0;
    hbm_apb_pslverr_1 = 'b0;

    hbm_apb_paddr_0   = 'b0;
    hbm_apb_pprot_0   = 'b0;
    hbm_apb_psel_0    = 'b0;
    hbm_apb_penable_0 = 'b0;
    hbm_apb_pwrite_0  = 'b0;
    hbm_apb_pwdata_0  = 'b0;
    hbm_apb_pstrb_0   = 'b0;
    hbm_apb_pready_0  = 'b0;
    hbm_apb_prdata_0  = 'b0;
    hbm_apb_pslverr_0 = 'b0;
  end

//=============================================================================
// C2C IO
//=============================================================================

  always_comb begin
    PCIE_EP_TXP    = 'b0;
    PCIE_EP_TXN    = 'b0;

    PCIE_RP_PERSTN = 'b0;
    PCIE_RP_TXP    = 'b0;
    PCIE_RP_TXN    = 'b0;
  end

endmodule // prospero
