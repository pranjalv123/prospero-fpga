
    module circuit#(
        parameter WIDTH = 32,        // Total width of the operand
        parameter FRAC_BITS = 16     // Number of fractional bits
    )(
        input logic clk,
        input logic reset,
        input logic [WIDTH-1:0] x,
        input logic [WIDTH-1:0] y,
        output logic [WIDTH-1:0] out
    );
    
        logic [WIDTH-1:0] out_0;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.95)
        ) inst_0 (
            .outp(out_0)
        );
        

        logic [WIDTH-1:0] out_1;
        assign out_1 = x;
        

        logic [WIDTH-1:0] out_2;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.13008)
        ) inst_2 (
            .outp(out_2)
        );
        

        logic [WIDTH-1:0] out_3;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3 (
            .a(out_1),
            .b(out_2),
            .outp(out_3)
        );        
        

        logic [WIDTH-1:0] out_4;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4 (
            .a(out_0),
            .b(out_3),
            .outp(out_4)
        );        
        

        logic [WIDTH-1:0] out_5;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.675)
        ) inst_5 (
            .outp(out_5)
        );
        

        logic [WIDTH-1:0] out_6;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6 (
            .a(out_5),
            .b(out_3),
            .outp(out_6)
        );        
        

        logic [WIDTH-1:0] out_7;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7 (
            .in(out_6),
            .outp(out_7)
        );
        

        logic [WIDTH-1:0] out_8;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_8 (
            .a(out_4),
            .b(out_7),
            .outp(out_8)
        );        
        

        logic [WIDTH-1:0] out_9;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.175)
        ) inst_9 (
            .outp(out_9)
        );
        

        logic [WIDTH-1:0] out_10;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_10 (
            .in(out_4),
            .outp(out_10)
        );
        

        logic [WIDTH-1:0] out_11;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_11 (
            .in(out_10),
            .outp(out_11)
        );
        

        logic [WIDTH-1:0] out_12;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.025)
        ) inst_12 (
            .outp(out_12)
        );
        

        logic [WIDTH-1:0] out_13;
        assign out_13 = y;
        

        logic [WIDTH-1:0] out_14;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_14 (
            .a(out_13),
            .b(out_2),
            .outp(out_14)
        );        
        

        logic [WIDTH-1:0] out_15;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_15 (
            .a(out_12),
            .b(out_14),
            .outp(out_15)
        );        
        

        logic [WIDTH-1:0] out_16;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_16 (
            .in(out_15),
            .outp(out_16)
        );
        

        logic [WIDTH-1:0] out_17;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_17 (
            .a(out_11),
            .b(out_16),
            .outp(out_17)
        );        
        

        logic [WIDTH-1:0] out_18;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_18 (
            .in(out_17),
            .outp(out_18)
        );
        

        logic [WIDTH-1:0] out_19;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_19 (
            .a(out_9),
            .b(out_18),
            .outp(out_19)
        );        
        

        logic [WIDTH-1:0] out_20;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_20 (
            .a(out_8),
            .b(out_19),
            .outp(out_20)
        );        
        

        logic [WIDTH-1:0] out_21;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.275)
        ) inst_21 (
            .outp(out_21)
        );
        

        logic [WIDTH-1:0] out_22;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_22 (
            .a(out_18),
            .b(out_21),
            .outp(out_22)
        );        
        

        logic [WIDTH-1:0] out_23;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_23 (
            .a(out_20),
            .b(out_22),
            .outp(out_23)
        );        
        

        logic [WIDTH-1:0] out_24;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.3)
        ) inst_24 (
            .outp(out_24)
        );
        

        logic [WIDTH-1:0] out_25;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_25 (
            .a(out_24),
            .b(out_14),
            .outp(out_25)
        );        
        

        logic [WIDTH-1:0] out_26;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_26 (
            .a(out_23),
            .b(out_25),
            .outp(out_26)
        );        
        

        logic [WIDTH-1:0] out_27;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.3)
        ) inst_27 (
            .outp(out_27)
        );
        

        logic [WIDTH-1:0] out_28;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_28 (
            .a(out_27),
            .b(out_14),
            .outp(out_28)
        );        
        

        logic [WIDTH-1:0] out_29;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_29 (
            .in(out_28),
            .outp(out_29)
        );
        

        logic [WIDTH-1:0] out_30;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_30 (
            .a(out_26),
            .b(out_29),
            .outp(out_30)
        );        
        

        logic [WIDTH-1:0] out_31;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.025)
        ) inst_31 (
            .outp(out_31)
        );
        

        logic [WIDTH-1:0] out_32;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_32 (
            .a(out_31),
            .b(out_3),
            .outp(out_32)
        );        
        

        logic [WIDTH-1:0] out_33;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.125)
        ) inst_33 (
            .outp(out_33)
        );
        

        logic [WIDTH-1:0] out_34;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_34 (
            .a(out_33),
            .b(out_3),
            .outp(out_34)
        );        
        

        logic [WIDTH-1:0] out_35;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_35 (
            .in(out_34),
            .outp(out_35)
        );
        

        logic [WIDTH-1:0] out_36;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_36 (
            .a(out_32),
            .b(out_35),
            .outp(out_36)
        );        
        

        logic [WIDTH-1:0] out_37;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_37 (
            .a(out_36),
            .b(out_25),
            .outp(out_37)
        );        
        

        logic [WIDTH-1:0] out_38;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_38 (
            .a(out_37),
            .b(out_29),
            .outp(out_38)
        );        
        

        logic [WIDTH-1:0] out_39;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_39 (
            .a(out_30),
            .b(out_38),
            .outp(out_39)
        );        
        

        logic [WIDTH-1:0] out_40;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.275)
        ) inst_40 (
            .outp(out_40)
        );
        

        logic [WIDTH-1:0] out_41;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_41 (
            .a(out_40),
            .b(out_3),
            .outp(out_41)
        );        
        

        logic [WIDTH-1:0] out_42;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.375)
        ) inst_42 (
            .outp(out_42)
        );
        

        logic [WIDTH-1:0] out_43;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_43 (
            .a(out_42),
            .b(out_3),
            .outp(out_43)
        );        
        

        logic [WIDTH-1:0] out_44;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_44 (
            .in(out_43),
            .outp(out_44)
        );
        

        logic [WIDTH-1:0] out_45;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_45 (
            .a(out_41),
            .b(out_44),
            .outp(out_45)
        );        
        

        logic [WIDTH-1:0] out_46;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_46 (
            .a(out_45),
            .b(out_25),
            .outp(out_46)
        );        
        

        logic [WIDTH-1:0] out_47;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_47 (
            .a(out_46),
            .b(out_29),
            .outp(out_47)
        );        
        

        logic [WIDTH-1:0] out_48;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_48 (
            .a(out_39),
            .b(out_47),
            .outp(out_48)
        );        
        

        logic [WIDTH-1:0] out_49;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.5)
        ) inst_49 (
            .outp(out_49)
        );
        

        logic [WIDTH-1:0] out_50;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_50 (
            .a(out_49),
            .b(out_14),
            .outp(out_50)
        );        
        

        logic [WIDTH-1:0] out_51;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.75)
        ) inst_51 (
            .outp(out_51)
        );
        

        logic [WIDTH-1:0] out_52;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_52 (
            .a(out_51),
            .b(out_14),
            .outp(out_52)
        );        
        

        logic [WIDTH-1:0] out_53;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_53 (
            .in(out_52),
            .outp(out_53)
        );
        

        logic [WIDTH-1:0] out_54;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_54 (
            .a(out_50),
            .b(out_53),
            .outp(out_54)
        );        
        

        logic [WIDTH-1:0] out_55;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5)
        ) inst_55 (
            .outp(out_55)
        );
        

        logic [WIDTH-1:0] out_56;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_56 (
            .a(out_55),
            .b(out_3),
            .outp(out_56)
        );        
        

        logic [WIDTH-1:0] out_57;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_57 (
            .a(out_54),
            .b(out_56),
            .outp(out_57)
        );        
        

        logic [WIDTH-1:0] out_58;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.6)
        ) inst_58 (
            .outp(out_58)
        );
        

        logic [WIDTH-1:0] out_59;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_59 (
            .a(out_58),
            .b(out_3),
            .outp(out_59)
        );        
        

        logic [WIDTH-1:0] out_60;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_60 (
            .in(out_59),
            .outp(out_60)
        );
        

        logic [WIDTH-1:0] out_61;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_61 (
            .a(out_57),
            .b(out_60),
            .outp(out_61)
        );        
        

        logic [WIDTH-1:0] out_62;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_62 (
            .a(out_48),
            .b(out_61),
            .outp(out_62)
        );        
        

        logic [WIDTH-1:0] out_63;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.4)
        ) inst_63 (
            .outp(out_63)
        );
        

        logic [WIDTH-1:0] out_64;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_64 (
            .a(out_63),
            .b(out_14),
            .outp(out_64)
        );        
        

        logic [WIDTH-1:0] out_65;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_65 (
            .in(out_64),
            .outp(out_65)
        );
        

        logic [WIDTH-1:0] out_66;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.7)
        ) inst_66 (
            .outp(out_66)
        );
        

        logic [WIDTH-1:0] out_67;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_67 (
            .a(out_66),
            .b(out_3),
            .outp(out_67)
        );        
        

        logic [WIDTH-1:0] out_68;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_68 (
            .a(out_65),
            .b(out_67),
            .outp(out_68)
        );        
        

        logic [WIDTH-1:0] out_69;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.2)
        ) inst_69 (
            .outp(out_69)
        );
        

        logic [WIDTH-1:0] out_70;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_70 (
            .a(out_69),
            .b(out_3),
            .outp(out_70)
        );        
        

        logic [WIDTH-1:0] out_71;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_71 (
            .in(out_70),
            .outp(out_71)
        );
        

        logic [WIDTH-1:0] out_72;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_72 (
            .a(out_68),
            .b(out_71),
            .outp(out_72)
        );        
        

        logic [WIDTH-1:0] out_73;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_73 (
            .a(out_72),
            .b(out_25),
            .outp(out_73)
        );        
        

        logic [WIDTH-1:0] out_74;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_74 (
            .a(out_62),
            .b(out_73),
            .outp(out_74)
        );        
        

        logic [WIDTH-1:0] out_75;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_75 (
            .a(out_67),
            .b(out_71),
            .outp(out_75)
        );        
        

        logic [WIDTH-1:0] out_76;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.2)
        ) inst_76 (
            .outp(out_76)
        );
        

        logic [WIDTH-1:0] out_77;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_77 (
            .a(out_76),
            .b(out_14),
            .outp(out_77)
        );        
        

        logic [WIDTH-1:0] out_78;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_78 (
            .a(out_75),
            .b(out_77),
            .outp(out_78)
        );        
        

        logic [WIDTH-1:0] out_79;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_79 (
            .a(out_78),
            .b(out_29),
            .outp(out_79)
        );        
        

        logic [WIDTH-1:0] out_80;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_80 (
            .a(out_74),
            .b(out_79),
            .outp(out_80)
        );        
        

        logic [WIDTH-1:0] out_81;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.9)
        ) inst_81 (
            .outp(out_81)
        );
        

        logic [WIDTH-1:0] out_82;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_82 (
            .a(out_81),
            .b(out_3),
            .outp(out_82)
        );        
        

        logic [WIDTH-1:0] out_83;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.0)
        ) inst_83 (
            .outp(out_83)
        );
        

        logic [WIDTH-1:0] out_84;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_84 (
            .a(out_83),
            .b(out_3),
            .outp(out_84)
        );        
        

        logic [WIDTH-1:0] out_85;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_85 (
            .in(out_84),
            .outp(out_85)
        );
        

        logic [WIDTH-1:0] out_86;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_86 (
            .a(out_82),
            .b(out_85),
            .outp(out_86)
        );        
        

        logic [WIDTH-1:0] out_87;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_87 (
            .a(out_86),
            .b(out_25),
            .outp(out_87)
        );        
        

        logic [WIDTH-1:0] out_88;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_88 (
            .a(out_87),
            .b(out_29),
            .outp(out_88)
        );        
        

        logic [WIDTH-1:0] out_89;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_89 (
            .a(out_80),
            .b(out_88),
            .outp(out_89)
        );        
        

        logic [WIDTH-1:0] out_90;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.2)
        ) inst_90 (
            .outp(out_90)
        );
        

        logic [WIDTH-1:0] out_91;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_91 (
            .a(out_90),
            .b(out_14),
            .outp(out_91)
        );        
        

        logic [WIDTH-1:0] out_92;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.2)
        ) inst_92 (
            .outp(out_92)
        );
        

        logic [WIDTH-1:0] out_93;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_93 (
            .a(out_92),
            .b(out_14),
            .outp(out_93)
        );        
        

        logic [WIDTH-1:0] out_94;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_94 (
            .in(out_93),
            .outp(out_94)
        );
        

        logic [WIDTH-1:0] out_95;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_95 (
            .a(out_91),
            .b(out_94),
            .outp(out_95)
        );        
        

        logic [WIDTH-1:0] out_96;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.7205)
        ) inst_96 (
            .outp(out_96)
        );
        

        logic [WIDTH-1:0] out_97;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_97 (
            .a(out_96),
            .b(out_3),
            .outp(out_97)
        );        
        

        logic [WIDTH-1:0] out_98;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_98 (
            .a(out_95),
            .b(out_97),
            .outp(out_98)
        );        
        

        logic [WIDTH-1:0] out_99;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.8205)
        ) inst_99 (
            .outp(out_99)
        );
        

        logic [WIDTH-1:0] out_100;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_100 (
            .a(out_3),
            .b(out_99),
            .outp(out_100)
        );        
        

        logic [WIDTH-1:0] out_101;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_101 (
            .a(out_98),
            .b(out_100),
            .outp(out_101)
        );        
        

        logic [WIDTH-1:0] out_102;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_102 (
            .a(out_89),
            .b(out_101),
            .outp(out_102)
        );        
        

        logic [WIDTH-1:0] out_103;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.65)
        ) inst_103 (
            .outp(out_103)
        );
        

        logic [WIDTH-1:0] out_104;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_104 (
            .a(out_103),
            .b(out_14),
            .outp(out_104)
        );        
        

        logic [WIDTH-1:0] out_105;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.75)
        ) inst_105 (
            .outp(out_105)
        );
        

        logic [WIDTH-1:0] out_106;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_106 (
            .a(out_105),
            .b(out_14),
            .outp(out_106)
        );        
        

        logic [WIDTH-1:0] out_107;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_107 (
            .in(out_106),
            .outp(out_107)
        );
        

        logic [WIDTH-1:0] out_108;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_108 (
            .a(out_104),
            .b(out_107),
            .outp(out_108)
        );        
        

        logic [WIDTH-1:0] out_109;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.54551)
        ) inst_109 (
            .outp(out_109)
        );
        

        logic [WIDTH-1:0] out_110;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_110 (
            .a(out_109),
            .b(out_3),
            .outp(out_110)
        );        
        

        logic [WIDTH-1:0] out_111;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_111 (
            .a(out_108),
            .b(out_110),
            .outp(out_111)
        );        
        

        logic [WIDTH-1:0] out_112;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.7205)
        ) inst_112 (
            .outp(out_112)
        );
        

        logic [WIDTH-1:0] out_113;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_113 (
            .a(out_3),
            .b(out_112),
            .outp(out_113)
        );        
        

        logic [WIDTH-1:0] out_114;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_114 (
            .a(out_111),
            .b(out_113),
            .outp(out_114)
        );        
        

        logic [WIDTH-1:0] out_115;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_115 (
            .a(out_102),
            .b(out_114),
            .outp(out_115)
        );        
        

        logic [WIDTH-1:0] out_116;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_116 (
            .a(out_94),
            .b(out_110),
            .outp(out_116)
        );        
        

        logic [WIDTH-1:0] out_117;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_117 (
            .a(out_116),
            .b(out_113),
            .outp(out_117)
        );        
        

        logic [WIDTH-1:0] out_118;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.1)
        ) inst_118 (
            .outp(out_118)
        );
        

        logic [WIDTH-1:0] out_119;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_119 (
            .a(out_118),
            .b(out_14),
            .outp(out_119)
        );        
        

        logic [WIDTH-1:0] out_120;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_120 (
            .a(out_117),
            .b(out_119),
            .outp(out_120)
        );        
        

        logic [WIDTH-1:0] out_121;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_121 (
            .a(out_115),
            .b(out_120),
            .outp(out_121)
        );        
        

        logic [WIDTH-1:0] out_122;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.53565)
        ) inst_122 (
            .outp(out_122)
        );
        

        logic [WIDTH-1:0] out_123;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.84553)
        ) inst_123 (
            .outp(out_123)
        );
        

        logic [WIDTH-1:0] out_124;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_124 (
            .a(out_13),
            .b(out_123),
            .outp(out_124)
        );        
        

        logic [WIDTH-1:0] out_125;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_125 (
            .a(out_122),
            .b(out_124),
            .outp(out_125)
        );        
        

        logic [WIDTH-1:0] out_126;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.47154)
        ) inst_126 (
            .outp(out_126)
        );
        

        logic [WIDTH-1:0] out_127;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_127 (
            .a(out_1),
            .b(out_126),
            .outp(out_127)
        );        
        

        logic [WIDTH-1:0] out_128;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_128 (
            .a(out_125),
            .b(out_127),
            .outp(out_128)
        );        
        

        logic [WIDTH-1:0] out_129;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.90565)
        ) inst_129 (
            .outp(out_129)
        );
        

        logic [WIDTH-1:0] out_130;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.03252)
        ) inst_130 (
            .outp(out_130)
        );
        

        logic [WIDTH-1:0] out_131;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_131 (
            .a(out_13),
            .b(out_130),
            .outp(out_131)
        );        
        

        logic [WIDTH-1:0] out_132;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_132 (
            .a(out_129),
            .b(out_131),
            .outp(out_132)
        );        
        

        logic [WIDTH-1:0] out_133;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_133 (
            .a(out_127),
            .b(out_132),
            .outp(out_133)
        );        
        

        logic [WIDTH-1:0] out_134;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_134 (
            .a(out_128),
            .b(out_133),
            .outp(out_134)
        );        
        

        logic [WIDTH-1:0] out_135;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.575)
        ) inst_135 (
            .outp(out_135)
        );
        

        logic [WIDTH-1:0] out_136;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.813008)
        ) inst_136 (
            .outp(out_136)
        );
        

        logic [WIDTH-1:0] out_137;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_137 (
            .a(out_13),
            .b(out_136),
            .outp(out_137)
        );        
        

        logic [WIDTH-1:0] out_138;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_138 (
            .a(out_135),
            .b(out_137),
            .outp(out_138)
        );        
        

        logic [WIDTH-1:0] out_139;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_139 (
            .in(out_138),
            .outp(out_139)
        );
        

        logic [WIDTH-1:0] out_140;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_140 (
            .a(out_134),
            .b(out_139),
            .outp(out_140)
        );        
        

        logic [WIDTH-1:0] out_141;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_141 (
            .a(out_121),
            .b(out_140),
            .outp(out_141)
        );        
        

        logic [WIDTH-1:0] out_142;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.24435)
        ) inst_142 (
            .outp(out_142)
        );
        

        logic [WIDTH-1:0] out_143;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_143 (
            .a(out_131),
            .b(out_142),
            .outp(out_143)
        );        
        

        logic [WIDTH-1:0] out_144;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_144 (
            .a(out_143),
            .b(out_127),
            .outp(out_144)
        );        
        

        logic [WIDTH-1:0] out_145;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_145 (
            .in(out_144),
            .outp(out_145)
        );
        

        logic [WIDTH-1:0] out_146;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.81935)
        ) inst_146 (
            .outp(out_146)
        );
        

        logic [WIDTH-1:0] out_147;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_147 (
            .a(out_146),
            .b(out_124),
            .outp(out_147)
        );        
        

        logic [WIDTH-1:0] out_148;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_148 (
            .a(out_147),
            .b(out_127),
            .outp(out_148)
        );        
        

        logic [WIDTH-1:0] out_149;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_149 (
            .a(out_145),
            .b(out_148),
            .outp(out_149)
        );        
        

        logic [WIDTH-1:0] out_150;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.63)
        ) inst_150 (
            .outp(out_150)
        );
        

        logic [WIDTH-1:0] out_151;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.813008)
        ) inst_151 (
            .outp(out_151)
        );
        

        logic [WIDTH-1:0] out_152;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_152 (
            .a(out_13),
            .b(out_151),
            .outp(out_152)
        );        
        

        logic [WIDTH-1:0] out_153;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_153 (
            .a(out_150),
            .b(out_152),
            .outp(out_153)
        );        
        

        logic [WIDTH-1:0] out_154;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_154 (
            .in(out_153),
            .outp(out_154)
        );
        

        logic [WIDTH-1:0] out_155;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_155 (
            .a(out_149),
            .b(out_154),
            .outp(out_155)
        );        
        

        logic [WIDTH-1:0] out_156;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_156 (
            .a(out_141),
            .b(out_155),
            .outp(out_156)
        );        
        

        logic [WIDTH-1:0] out_157;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.81935)
        ) inst_157 (
            .outp(out_157)
        );
        

        logic [WIDTH-1:0] out_158;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_158 (
            .a(out_157),
            .b(out_124),
            .outp(out_158)
        );        
        

        logic [WIDTH-1:0] out_159;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_159 (
            .a(out_158),
            .b(out_127),
            .outp(out_159)
        );        
        

        logic [WIDTH-1:0] out_160;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_160 (
            .in(out_159),
            .outp(out_160)
        );
        

        logic [WIDTH-1:0] out_161;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_161 (
            .a(out_144),
            .b(out_160),
            .outp(out_161)
        );        
        

        logic [WIDTH-1:0] out_162;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_162 (
            .a(out_161),
            .b(out_153),
            .outp(out_162)
        );        
        

        logic [WIDTH-1:0] out_163;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_163 (
            .a(out_156),
            .b(out_162),
            .outp(out_163)
        );        
        

        logic [WIDTH-1:0] out_164;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.18935)
        ) inst_164 (
            .outp(out_164)
        );
        

        logic [WIDTH-1:0] out_165;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_165 (
            .a(out_131),
            .b(out_164),
            .outp(out_165)
        );        
        

        logic [WIDTH-1:0] out_166;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_166 (
            .a(out_165),
            .b(out_127),
            .outp(out_166)
        );        
        

        logic [WIDTH-1:0] out_167;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_167 (
            .a(out_160),
            .b(out_166),
            .outp(out_167)
        );        
        

        logic [WIDTH-1:0] out_168;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_168 (
            .a(out_167),
            .b(out_138),
            .outp(out_168)
        );        
        

        logic [WIDTH-1:0] out_169;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_169 (
            .a(out_163),
            .b(out_168),
            .outp(out_169)
        );        
        

        logic [WIDTH-1:0] out_170;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_170 (
            .in(out_166),
            .outp(out_170)
        );
        

        logic [WIDTH-1:0] out_171;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_171 (
            .a(out_148),
            .b(out_170),
            .outp(out_171)
        );        
        

        logic [WIDTH-1:0] out_172;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_172 (
            .a(out_171),
            .b(out_139),
            .outp(out_172)
        );        
        

        logic [WIDTH-1:0] out_173;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_173 (
            .a(out_169),
            .b(out_172),
            .outp(out_173)
        );        
        

        logic [WIDTH-1:0] out_174;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.842)
        ) inst_174 (
            .outp(out_174)
        );
        

        logic [WIDTH-1:0] out_175;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_175 (
            .a(out_174),
            .b(out_3),
            .outp(out_175)
        );        
        

        logic [WIDTH-1:0] out_176;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_176 (
            .in(out_175),
            .outp(out_176)
        );
        

        logic [WIDTH-1:0] out_177;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_177 (
            .a(out_176),
            .b(out_16),
            .outp(out_177)
        );        
        

        logic [WIDTH-1:0] out_178;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_178 (
            .in(out_177),
            .outp(out_178)
        );
        

        logic [WIDTH-1:0] out_179;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_179 (
            .a(out_9),
            .b(out_178),
            .outp(out_179)
        );        
        

        logic [WIDTH-1:0] out_180;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_180 (
            .a(out_178),
            .b(out_21),
            .outp(out_180)
        );        
        

        logic [WIDTH-1:0] out_181;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_181 (
            .a(out_179),
            .b(out_180),
            .outp(out_181)
        );        
        

        logic [WIDTH-1:0] out_182;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_182 (
            .a(out_173),
            .b(out_181),
            .outp(out_182)
        );        
        

        logic [WIDTH-1:0] out_183;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.475)
        ) inst_183 (
            .outp(out_183)
        );
        

        logic [WIDTH-1:0] out_184;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_184 (
            .a(out_183),
            .b(out_3),
            .outp(out_184)
        );        
        

        logic [WIDTH-1:0] out_185;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.575)
        ) inst_185 (
            .outp(out_185)
        );
        

        logic [WIDTH-1:0] out_186;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_186 (
            .a(out_185),
            .b(out_3),
            .outp(out_186)
        );        
        

        logic [WIDTH-1:0] out_187;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_187 (
            .in(out_186),
            .outp(out_187)
        );
        

        logic [WIDTH-1:0] out_188;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_188 (
            .a(out_184),
            .b(out_187),
            .outp(out_188)
        );        
        

        logic [WIDTH-1:0] out_189;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_189 (
            .a(out_188),
            .b(out_52),
            .outp(out_189)
        );        
        

        logic [WIDTH-1:0] out_190;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_190 (
            .a(out_189),
            .b(out_29),
            .outp(out_190)
        );        
        

        logic [WIDTH-1:0] out_191;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_191 (
            .a(out_182),
            .b(out_190),
            .outp(out_191)
        );        
        

        logic [WIDTH-1:0] out_192;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.12857)
        ) inst_192 (
            .outp(out_192)
        );
        

        logic [WIDTH-1:0] out_193;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(11.6144)
        ) inst_193 (
            .outp(out_193)
        );
        

        logic [WIDTH-1:0] out_194;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_194 (
            .a(out_1),
            .b(out_193),
            .outp(out_194)
        );        
        

        logic [WIDTH-1:0] out_195;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_195 (
            .a(out_192),
            .b(out_194),
            .outp(out_195)
        );        
        

        logic [WIDTH-1:0] out_196;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.67857)
        ) inst_196 (
            .outp(out_196)
        );
        

        logic [WIDTH-1:0] out_197;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_197 (
            .a(out_196),
            .b(out_194),
            .outp(out_197)
        );        
        

        logic [WIDTH-1:0] out_198;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_198 (
            .in(out_197),
            .outp(out_198)
        );
        

        logic [WIDTH-1:0] out_199;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_199 (
            .a(out_195),
            .b(out_198),
            .outp(out_199)
        );        
        

        logic [WIDTH-1:0] out_200;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.45)
        ) inst_200 (
            .outp(out_200)
        );
        

        logic [WIDTH-1:0] out_201;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_201 (
            .in(out_28),
            .outp(out_201)
        );
        

        logic [WIDTH-1:0] out_202;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.91072)
        ) inst_202 (
            .outp(out_202)
        );
        

        logic [WIDTH-1:0] out_203;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(14.518)
        ) inst_203 (
            .outp(out_203)
        );
        

        logic [WIDTH-1:0] out_204;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_204 (
            .a(out_1),
            .b(out_203),
            .outp(out_204)
        );        
        

        logic [WIDTH-1:0] out_205;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_205 (
            .a(out_202),
            .b(out_204),
            .outp(out_205)
        );        
        

        logic [WIDTH-1:0] out_206;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_206 (
            .in(out_205),
            .outp(out_206)
        );
        

        logic [WIDTH-1:0] out_207;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_207 (
            .a(out_201),
            .b(out_206),
            .outp(out_207)
        );        
        

        logic [WIDTH-1:0] out_208;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_208 (
            .in(out_207),
            .outp(out_208)
        );
        

        logic [WIDTH-1:0] out_209;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_209 (
            .a(out_200),
            .b(out_208),
            .outp(out_209)
        );        
        

        logic [WIDTH-1:0] out_210;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_210 (
            .a(out_199),
            .b(out_209),
            .outp(out_210)
        );        
        

        logic [WIDTH-1:0] out_211;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_211 (
            .in(out_195),
            .outp(out_211)
        );
        

        logic [WIDTH-1:0] out_212;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_212 (
            .a(out_201),
            .b(out_211),
            .outp(out_212)
        );        
        

        logic [WIDTH-1:0] out_213;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_213 (
            .in(out_212),
            .outp(out_213)
        );
        

        logic [WIDTH-1:0] out_214;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.55)
        ) inst_214 (
            .outp(out_214)
        );
        

        logic [WIDTH-1:0] out_215;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_215 (
            .a(out_213),
            .b(out_214),
            .outp(out_215)
        );        
        

        logic [WIDTH-1:0] out_216;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_216 (
            .a(out_210),
            .b(out_215),
            .outp(out_216)
        );        
        

        logic [WIDTH-1:0] out_217;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_217 (
            .a(out_216),
            .b(out_52),
            .outp(out_217)
        );        
        

        logic [WIDTH-1:0] out_218;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_218 (
            .a(out_217),
            .b(out_29),
            .outp(out_218)
        );        
        

        logic [WIDTH-1:0] out_219;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_219 (
            .a(out_191),
            .b(out_218),
            .outp(out_219)
        );        
        

        logic [WIDTH-1:0] out_220;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.775)
        ) inst_220 (
            .outp(out_220)
        );
        

        logic [WIDTH-1:0] out_221;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_221 (
            .a(out_220),
            .b(out_3),
            .outp(out_221)
        );        
        

        logic [WIDTH-1:0] out_222;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_222 (
            .in(out_221),
            .outp(out_222)
        );
        

        logic [WIDTH-1:0] out_223;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.675)
        ) inst_223 (
            .outp(out_223)
        );
        

        logic [WIDTH-1:0] out_224;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_224 (
            .a(out_223),
            .b(out_3),
            .outp(out_224)
        );        
        

        logic [WIDTH-1:0] out_225;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_225 (
            .a(out_222),
            .b(out_224),
            .outp(out_225)
        );        
        

        logic [WIDTH-1:0] out_226;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_226 (
            .a(out_225),
            .b(out_25),
            .outp(out_226)
        );        
        

        logic [WIDTH-1:0] out_227;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_227 (
            .a(out_226),
            .b(out_29),
            .outp(out_227)
        );        
        

        logic [WIDTH-1:0] out_228;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_228 (
            .a(out_219),
            .b(out_227),
            .outp(out_228)
        );        
        

        logic [WIDTH-1:0] out_229;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_229 (
            .a(out_221),
            .b(out_10),
            .outp(out_229)
        );        
        

        logic [WIDTH-1:0] out_230;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_230 (
            .a(out_229),
            .b(out_52),
            .outp(out_230)
        );        
        

        logic [WIDTH-1:0] out_231;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.85)
        ) inst_231 (
            .outp(out_231)
        );
        

        logic [WIDTH-1:0] out_232;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_232 (
            .a(out_231),
            .b(out_14),
            .outp(out_232)
        );        
        

        logic [WIDTH-1:0] out_233;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_233 (
            .in(out_232),
            .outp(out_233)
        );
        

        logic [WIDTH-1:0] out_234;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_234 (
            .a(out_230),
            .b(out_233),
            .outp(out_234)
        );        
        

        logic [WIDTH-1:0] out_235;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_235 (
            .a(out_228),
            .b(out_234),
            .outp(out_235)
        );        
        

        logic [WIDTH-1:0] out_236;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_236 (
            .a(out_229),
            .b(out_77),
            .outp(out_236)
        );        
        

        logic [WIDTH-1:0] out_237;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_237 (
            .a(out_236),
            .b(out_29),
            .outp(out_237)
        );        
        

        logic [WIDTH-1:0] out_238;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_238 (
            .a(out_235),
            .b(out_237),
            .outp(out_238)
        );        
        

        logic [WIDTH-1:0] out_239;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.33245)
        ) inst_239 (
            .outp(out_239)
        );
        

        logic [WIDTH-1:0] out_240;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.61337)
        ) inst_240 (
            .outp(out_240)
        );
        

        logic [WIDTH-1:0] out_241;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_241 (
            .a(out_1),
            .b(out_240),
            .outp(out_241)
        );        
        

        logic [WIDTH-1:0] out_242;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_242 (
            .a(out_239),
            .b(out_241),
            .outp(out_242)
        );        
        

        logic [WIDTH-1:0] out_243;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_243 (
            .in(out_242),
            .outp(out_243)
        );
        

        logic [WIDTH-1:0] out_244;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.815)
        ) inst_244 (
            .outp(out_244)
        );
        

        logic [WIDTH-1:0] out_245;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_245 (
            .a(out_244),
            .b(out_14),
            .outp(out_245)
        );        
        

        logic [WIDTH-1:0] out_246;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_246 (
            .in(out_245),
            .outp(out_246)
        );
        

        logic [WIDTH-1:0] out_247;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_247 (
            .in(out_246),
            .outp(out_247)
        );
        

        logic [WIDTH-1:0] out_248;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_248 (
            .a(out_243),
            .b(out_247),
            .outp(out_248)
        );        
        

        logic [WIDTH-1:0] out_249;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_249 (
            .in(out_248),
            .outp(out_249)
        );
        

        logic [WIDTH-1:0] out_250;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0625)
        ) inst_250 (
            .outp(out_250)
        );
        

        logic [WIDTH-1:0] out_251;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_251 (
            .a(out_249),
            .b(out_250),
            .outp(out_251)
        );        
        

        logic [WIDTH-1:0] out_252;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.975)
        ) inst_252 (
            .outp(out_252)
        );
        

        logic [WIDTH-1:0] out_253;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_253 (
            .a(out_252),
            .b(out_14),
            .outp(out_253)
        );        
        

        logic [WIDTH-1:0] out_254;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_254 (
            .in(out_253),
            .outp(out_254)
        );
        

        logic [WIDTH-1:0] out_255;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.8125)
        ) inst_255 (
            .outp(out_255)
        );
        

        logic [WIDTH-1:0] out_256;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_256 (
            .a(out_255),
            .b(out_14),
            .outp(out_256)
        );        
        

        logic [WIDTH-1:0] out_257;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_257 (
            .a(out_254),
            .b(out_256),
            .outp(out_257)
        );        
        

        logic [WIDTH-1:0] out_258;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.00117)
        ) inst_258 (
            .outp(out_258)
        );
        

        logic [WIDTH-1:0] out_259;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.42005)
        ) inst_259 (
            .outp(out_259)
        );
        

        logic [WIDTH-1:0] out_260;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_260 (
            .a(out_1),
            .b(out_259),
            .outp(out_260)
        );        
        

        logic [WIDTH-1:0] out_261;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_261 (
            .a(out_258),
            .b(out_260),
            .outp(out_261)
        );        
        

        logic [WIDTH-1:0] out_262;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_262 (
            .a(out_257),
            .b(out_261),
            .outp(out_262)
        );        
        

        logic [WIDTH-1:0] out_263;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.16367)
        ) inst_263 (
            .outp(out_263)
        );
        

        logic [WIDTH-1:0] out_264;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_264 (
            .a(out_260),
            .b(out_263),
            .outp(out_264)
        );        
        

        logic [WIDTH-1:0] out_265;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_265 (
            .a(out_262),
            .b(out_264),
            .outp(out_265)
        );        
        

        logic [WIDTH-1:0] out_266;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_266 (
            .a(out_251),
            .b(out_265),
            .outp(out_266)
        );        
        

        logic [WIDTH-1:0] out_267;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_267 (
            .in(out_266),
            .outp(out_267)
        );
        

        logic [WIDTH-1:0] out_268;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.8125)
        ) inst_268 (
            .outp(out_268)
        );
        

        logic [WIDTH-1:0] out_269;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_269 (
            .a(out_268),
            .b(out_14),
            .outp(out_269)
        );        
        

        logic [WIDTH-1:0] out_270;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_270 (
            .in(out_269),
            .outp(out_270)
        );
        

        logic [WIDTH-1:0] out_271;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_271 (
            .in(out_270),
            .outp(out_271)
        );
        

        logic [WIDTH-1:0] out_272;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_272 (
            .in(out_261),
            .outp(out_272)
        );
        

        logic [WIDTH-1:0] out_273;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_273 (
            .a(out_271),
            .b(out_272),
            .outp(out_273)
        );        
        

        logic [WIDTH-1:0] out_274;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_274 (
            .in(out_273),
            .outp(out_274)
        );
        

        logic [WIDTH-1:0] out_275;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.1625)
        ) inst_275 (
            .outp(out_275)
        );
        

        logic [WIDTH-1:0] out_276;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_276 (
            .a(out_274),
            .b(out_275),
            .outp(out_276)
        );        
        

        logic [WIDTH-1:0] out_277;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_277 (
            .a(out_267),
            .b(out_276),
            .outp(out_277)
        );        
        

        logic [WIDTH-1:0] out_278;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_278 (
            .a(out_238),
            .b(out_277),
            .outp(out_278)
        );        
        

        logic [WIDTH-1:0] out_279;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.0375)
        ) inst_279 (
            .outp(out_279)
        );
        

        logic [WIDTH-1:0] out_280;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_280 (
            .a(out_279),
            .b(out_14),
            .outp(out_280)
        );        
        

        logic [WIDTH-1:0] out_281;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_281 (
            .in(out_280),
            .outp(out_281)
        );
        

        logic [WIDTH-1:0] out_282;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.00117)
        ) inst_282 (
            .outp(out_282)
        );
        

        logic [WIDTH-1:0] out_283;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_283 (
            .a(out_260),
            .b(out_282),
            .outp(out_283)
        );        
        

        logic [WIDTH-1:0] out_284;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_284 (
            .a(out_281),
            .b(out_283),
            .outp(out_284)
        );        
        

        logic [WIDTH-1:0] out_285;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.83867)
        ) inst_285 (
            .outp(out_285)
        );
        

        logic [WIDTH-1:0] out_286;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_286 (
            .a(out_285),
            .b(out_260),
            .outp(out_286)
        );        
        

        logic [WIDTH-1:0] out_287;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_287 (
            .a(out_284),
            .b(out_286),
            .outp(out_287)
        );        
        

        logic [WIDTH-1:0] out_288;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.875)
        ) inst_288 (
            .outp(out_288)
        );
        

        logic [WIDTH-1:0] out_289;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_289 (
            .a(out_288),
            .b(out_14),
            .outp(out_289)
        );        
        

        logic [WIDTH-1:0] out_290;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_290 (
            .a(out_287),
            .b(out_289),
            .outp(out_290)
        );        
        

        logic [WIDTH-1:0] out_291;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.035)
        ) inst_291 (
            .outp(out_291)
        );
        

        logic [WIDTH-1:0] out_292;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_292 (
            .a(out_291),
            .b(out_14),
            .outp(out_292)
        );        
        

        logic [WIDTH-1:0] out_293;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_293 (
            .in(out_292),
            .outp(out_293)
        );
        

        logic [WIDTH-1:0] out_294;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.33578)
        ) inst_294 (
            .outp(out_294)
        );
        

        logic [WIDTH-1:0] out_295;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_295 (
            .a(out_241),
            .b(out_294),
            .outp(out_295)
        );        
        

        logic [WIDTH-1:0] out_296;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_296 (
            .in(out_295),
            .outp(out_296)
        );
        

        logic [WIDTH-1:0] out_297;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_297 (
            .a(out_293),
            .b(out_296),
            .outp(out_297)
        );        
        

        logic [WIDTH-1:0] out_298;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_298 (
            .in(out_297),
            .outp(out_298)
        );
        

        logic [WIDTH-1:0] out_299;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_299 (
            .a(out_298),
            .b(out_250),
            .outp(out_299)
        );        
        

        logic [WIDTH-1:0] out_300;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_300 (
            .a(out_290),
            .b(out_299),
            .outp(out_300)
        );        
        

        logic [WIDTH-1:0] out_301;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_301 (
            .in(out_300),
            .outp(out_301)
        );
        

        logic [WIDTH-1:0] out_302;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.0375)
        ) inst_302 (
            .outp(out_302)
        );
        

        logic [WIDTH-1:0] out_303;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_303 (
            .a(out_302),
            .b(out_14),
            .outp(out_303)
        );        
        

        logic [WIDTH-1:0] out_304;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_304 (
            .in(out_303),
            .outp(out_304)
        );
        

        logic [WIDTH-1:0] out_305;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_305 (
            .in(out_283),
            .outp(out_305)
        );
        

        logic [WIDTH-1:0] out_306;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_306 (
            .a(out_304),
            .b(out_305),
            .outp(out_306)
        );        
        

        logic [WIDTH-1:0] out_307;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_307 (
            .in(out_306),
            .outp(out_307)
        );
        

        logic [WIDTH-1:0] out_308;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_308 (
            .a(out_307),
            .b(out_275),
            .outp(out_308)
        );        
        

        logic [WIDTH-1:0] out_309;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_309 (
            .a(out_301),
            .b(out_308),
            .outp(out_309)
        );        
        

        logic [WIDTH-1:0] out_310;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_310 (
            .a(out_278),
            .b(out_309),
            .outp(out_310)
        );        
        

        logic [WIDTH-1:0] out_311;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.95)
        ) inst_311 (
            .outp(out_311)
        );
        

        logic [WIDTH-1:0] out_312;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_312 (
            .a(out_311),
            .b(out_14),
            .outp(out_312)
        );        
        

        logic [WIDTH-1:0] out_313;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_313 (
            .in(out_312),
            .outp(out_313)
        );
        

        logic [WIDTH-1:0] out_314;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_314 (
            .a(out_91),
            .b(out_313),
            .outp(out_314)
        );        
        

        logic [WIDTH-1:0] out_315;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.808)
        ) inst_315 (
            .outp(out_315)
        );
        

        logic [WIDTH-1:0] out_316;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_316 (
            .a(out_3),
            .b(out_315),
            .outp(out_316)
        );        
        

        logic [WIDTH-1:0] out_317;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_317 (
            .a(out_314),
            .b(out_316),
            .outp(out_317)
        );        
        

        logic [WIDTH-1:0] out_318;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.708)
        ) inst_318 (
            .outp(out_318)
        );
        

        logic [WIDTH-1:0] out_319;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_319 (
            .a(out_318),
            .b(out_3),
            .outp(out_319)
        );        
        

        logic [WIDTH-1:0] out_320;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_320 (
            .a(out_317),
            .b(out_319),
            .outp(out_320)
        );        
        

        logic [WIDTH-1:0] out_321;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_321 (
            .a(out_310),
            .b(out_320),
            .outp(out_321)
        );        
        

        logic [WIDTH-1:0] out_322;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.55)
        ) inst_322 (
            .outp(out_322)
        );
        

        logic [WIDTH-1:0] out_323;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_323 (
            .a(out_322),
            .b(out_14),
            .outp(out_323)
        );        
        

        logic [WIDTH-1:0] out_324;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_324 (
            .in(out_104),
            .outp(out_324)
        );
        

        logic [WIDTH-1:0] out_325;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_325 (
            .a(out_323),
            .b(out_324),
            .outp(out_325)
        );        
        

        logic [WIDTH-1:0] out_326;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.958)
        ) inst_326 (
            .outp(out_326)
        );
        

        logic [WIDTH-1:0] out_327;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_327 (
            .a(out_3),
            .b(out_326),
            .outp(out_327)
        );        
        

        logic [WIDTH-1:0] out_328;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_328 (
            .a(out_325),
            .b(out_327),
            .outp(out_328)
        );        
        

        logic [WIDTH-1:0] out_329;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.558)
        ) inst_329 (
            .outp(out_329)
        );
        

        logic [WIDTH-1:0] out_330;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_330 (
            .a(out_329),
            .b(out_3),
            .outp(out_330)
        );        
        

        logic [WIDTH-1:0] out_331;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_331 (
            .a(out_328),
            .b(out_330),
            .outp(out_331)
        );        
        

        logic [WIDTH-1:0] out_332;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_332 (
            .a(out_321),
            .b(out_331),
            .outp(out_332)
        );        
        

        logic [WIDTH-1:0] out_333;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_333 (
            .a(out_94),
            .b(out_312),
            .outp(out_333)
        );        
        

        logic [WIDTH-1:0] out_334;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_334 (
            .a(out_333),
            .b(out_327),
            .outp(out_334)
        );        
        

        logic [WIDTH-1:0] out_335;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_335 (
            .a(out_334),
            .b(out_330),
            .outp(out_335)
        );        
        

        logic [WIDTH-1:0] out_336;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.15)
        ) inst_336 (
            .outp(out_336)
        );
        

        logic [WIDTH-1:0] out_337;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_337 (
            .in(out_312),
            .outp(out_337)
        );
        

        logic [WIDTH-1:0] out_338;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_338 (
            .in(out_327),
            .outp(out_338)
        );
        

        logic [WIDTH-1:0] out_339;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_339 (
            .a(out_337),
            .b(out_338),
            .outp(out_339)
        );        
        

        logic [WIDTH-1:0] out_340;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_340 (
            .in(out_339),
            .outp(out_340)
        );
        

        logic [WIDTH-1:0] out_341;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_341 (
            .a(out_336),
            .b(out_340),
            .outp(out_341)
        );        
        

        logic [WIDTH-1:0] out_342;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_342 (
            .a(out_335),
            .b(out_341),
            .outp(out_342)
        );        
        

        logic [WIDTH-1:0] out_343;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.25)
        ) inst_343 (
            .outp(out_343)
        );
        

        logic [WIDTH-1:0] out_344;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_344 (
            .a(out_340),
            .b(out_343),
            .outp(out_344)
        );        
        

        logic [WIDTH-1:0] out_345;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_345 (
            .a(out_342),
            .b(out_344),
            .outp(out_345)
        );        
        

        logic [WIDTH-1:0] out_346;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_346 (
            .a(out_332),
            .b(out_345),
            .outp(out_346)
        );        
        

        logic [WIDTH-1:0] out_347;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.8205)
        ) inst_347 (
            .outp(out_347)
        );
        

        logic [WIDTH-1:0] out_348;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_348 (
            .a(out_347),
            .b(out_3),
            .outp(out_348)
        );        
        

        logic [WIDTH-1:0] out_349;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_349 (
            .a(out_95),
            .b(out_348),
            .outp(out_349)
        );        
        

        logic [WIDTH-1:0] out_350;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.5455)
        ) inst_350 (
            .outp(out_350)
        );
        

        logic [WIDTH-1:0] out_351;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_351 (
            .a(out_3),
            .b(out_350),
            .outp(out_351)
        );        
        

        logic [WIDTH-1:0] out_352;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_352 (
            .a(out_349),
            .b(out_351),
            .outp(out_352)
        );        
        

        logic [WIDTH-1:0] out_353;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.925)
        ) inst_353 (
            .outp(out_353)
        );
        

        logic [WIDTH-1:0] out_354;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_354 (
            .a(out_353),
            .b(out_14),
            .outp(out_354)
        );        
        

        logic [WIDTH-1:0] out_355;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_355 (
            .in(out_354),
            .outp(out_355)
        );
        

        logic [WIDTH-1:0] out_356;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_356 (
            .in(out_110),
            .outp(out_356)
        );
        

        logic [WIDTH-1:0] out_357;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_357 (
            .a(out_355),
            .b(out_356),
            .outp(out_357)
        );        
        

        logic [WIDTH-1:0] out_358;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_358 (
            .in(out_357),
            .outp(out_358)
        );
        

        logic [WIDTH-1:0] out_359;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_359 (
            .a(out_9),
            .b(out_358),
            .outp(out_359)
        );        
        

        logic [WIDTH-1:0] out_360;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_360 (
            .a(out_352),
            .b(out_359),
            .outp(out_360)
        );        
        

        logic [WIDTH-1:0] out_361;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_361 (
            .a(out_358),
            .b(out_21),
            .outp(out_361)
        );        
        

        logic [WIDTH-1:0] out_362;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_362 (
            .a(out_360),
            .b(out_361),
            .outp(out_362)
        );        
        

        logic [WIDTH-1:0] out_363;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_363 (
            .a(out_346),
            .b(out_362),
            .outp(out_363)
        );        
        

        logic [WIDTH-1:0] out_364;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_364 (
            .a(out_94),
            .b(out_289),
            .outp(out_364)
        );        
        

        logic [WIDTH-1:0] out_365;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.1955)
        ) inst_365 (
            .outp(out_365)
        );
        

        logic [WIDTH-1:0] out_366;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_366 (
            .a(out_3),
            .b(out_365),
            .outp(out_366)
        );        
        

        logic [WIDTH-1:0] out_367;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_367 (
            .a(out_364),
            .b(out_366),
            .outp(out_367)
        );        
        

        logic [WIDTH-1:0] out_368;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.0955)
        ) inst_368 (
            .outp(out_368)
        );
        

        logic [WIDTH-1:0] out_369;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_369 (
            .a(out_368),
            .b(out_3),
            .outp(out_369)
        );        
        

        logic [WIDTH-1:0] out_370;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_370 (
            .a(out_367),
            .b(out_369),
            .outp(out_370)
        );        
        

        logic [WIDTH-1:0] out_371;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_371 (
            .a(out_363),
            .b(out_370),
            .outp(out_371)
        );        
        

        logic [WIDTH-1:0] out_372;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_372 (
            .a(out_94),
            .b(out_104),
            .outp(out_372)
        );        
        

        logic [WIDTH-1:0] out_373;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.7455)
        ) inst_373 (
            .outp(out_373)
        );
        

        logic [WIDTH-1:0] out_374;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_374 (
            .a(out_3),
            .b(out_373),
            .outp(out_374)
        );        
        

        logic [WIDTH-1:0] out_375;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_375 (
            .a(out_372),
            .b(out_374),
            .outp(out_375)
        );        
        

        logic [WIDTH-1:0] out_376;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.6455)
        ) inst_376 (
            .outp(out_376)
        );
        

        logic [WIDTH-1:0] out_377;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_377 (
            .a(out_376),
            .b(out_3),
            .outp(out_377)
        );        
        

        logic [WIDTH-1:0] out_378;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_378 (
            .a(out_375),
            .b(out_377),
            .outp(out_378)
        );        
        

        logic [WIDTH-1:0] out_379;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_379 (
            .a(out_371),
            .b(out_378),
            .outp(out_379)
        );        
        

        logic [WIDTH-1:0] out_380;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_380 (
            .a(out_104),
            .b(out_366),
            .outp(out_380)
        );        
        

        logic [WIDTH-1:0] out_381;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_381 (
            .a(out_380),
            .b(out_377),
            .outp(out_381)
        );        
        

        logic [WIDTH-1:0] out_382;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_382 (
            .in(out_289),
            .outp(out_382)
        );
        

        logic [WIDTH-1:0] out_383;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_383 (
            .a(out_381),
            .b(out_382),
            .outp(out_383)
        );        
        

        logic [WIDTH-1:0] out_384;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.9205)
        ) inst_384 (
            .outp(out_384)
        );
        

        logic [WIDTH-1:0] out_385;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_385 (
            .a(out_3),
            .b(out_384),
            .outp(out_385)
        );        
        

        logic [WIDTH-1:0] out_386;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_386 (
            .in(out_385),
            .outp(out_386)
        );
        

        logic [WIDTH-1:0] out_387;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_387 (
            .a(out_355),
            .b(out_386),
            .outp(out_387)
        );        
        

        logic [WIDTH-1:0] out_388;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_388 (
            .in(out_387),
            .outp(out_388)
        );
        

        logic [WIDTH-1:0] out_389;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_389 (
            .a(out_9),
            .b(out_388),
            .outp(out_389)
        );        
        

        logic [WIDTH-1:0] out_390;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_390 (
            .a(out_383),
            .b(out_389),
            .outp(out_390)
        );        
        

        logic [WIDTH-1:0] out_391;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_391 (
            .a(out_388),
            .b(out_21),
            .outp(out_391)
        );        
        

        logic [WIDTH-1:0] out_392;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_392 (
            .a(out_390),
            .b(out_391),
            .outp(out_392)
        );        
        

        logic [WIDTH-1:0] out_393;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_393 (
            .a(out_379),
            .b(out_392),
            .outp(out_393)
        );        
        

        logic [WIDTH-1:0] out_394;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5455)
        ) inst_394 (
            .outp(out_394)
        );
        

        logic [WIDTH-1:0] out_395;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_395 (
            .a(out_3),
            .b(out_394),
            .outp(out_395)
        );        
        

        logic [WIDTH-1:0] out_396;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_396 (
            .a(out_372),
            .b(out_395),
            .outp(out_396)
        );        
        

        logic [WIDTH-1:0] out_397;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.4455)
        ) inst_397 (
            .outp(out_397)
        );
        

        logic [WIDTH-1:0] out_398;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_398 (
            .a(out_397),
            .b(out_3),
            .outp(out_398)
        );        
        

        logic [WIDTH-1:0] out_399;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_399 (
            .a(out_396),
            .b(out_398),
            .outp(out_399)
        );        
        

        logic [WIDTH-1:0] out_400;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_400 (
            .a(out_393),
            .b(out_399),
            .outp(out_400)
        );        
        

        logic [WIDTH-1:0] out_401;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.925)
        ) inst_401 (
            .outp(out_401)
        );
        

        logic [WIDTH-1:0] out_402;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_402 (
            .a(out_401),
            .b(out_14),
            .outp(out_402)
        );        
        

        logic [WIDTH-1:0] out_403;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_403 (
            .in(out_402),
            .outp(out_403)
        );
        

        logic [WIDTH-1:0] out_404;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_404 (
            .a(out_104),
            .b(out_403),
            .outp(out_404)
        );        
        

        logic [WIDTH-1:0] out_405;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.0955)
        ) inst_405 (
            .outp(out_405)
        );
        

        logic [WIDTH-1:0] out_406;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_406 (
            .a(out_3),
            .b(out_405),
            .outp(out_406)
        );        
        

        logic [WIDTH-1:0] out_407;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_407 (
            .a(out_404),
            .b(out_406),
            .outp(out_407)
        );        
        

        logic [WIDTH-1:0] out_408;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.9955)
        ) inst_408 (
            .outp(out_408)
        );
        

        logic [WIDTH-1:0] out_409;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_409 (
            .a(out_408),
            .b(out_3),
            .outp(out_409)
        );        
        

        logic [WIDTH-1:0] out_410;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_410 (
            .a(out_407),
            .b(out_409),
            .outp(out_410)
        );        
        

        logic [WIDTH-1:0] out_411;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_411 (
            .a(out_400),
            .b(out_410),
            .outp(out_411)
        );        
        

        logic [WIDTH-1:0] out_412;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_412 (
            .a(out_94),
            .b(out_354),
            .outp(out_412)
        );        
        

        logic [WIDTH-1:0] out_413;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_413 (
            .a(out_412),
            .b(out_395),
            .outp(out_413)
        );        
        

        logic [WIDTH-1:0] out_414;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_414 (
            .a(out_413),
            .b(out_409),
            .outp(out_414)
        );        
        

        logic [WIDTH-1:0] out_415;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.2705)
        ) inst_415 (
            .outp(out_415)
        );
        

        logic [WIDTH-1:0] out_416;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_416 (
            .a(out_3),
            .b(out_415),
            .outp(out_416)
        );        
        

        logic [WIDTH-1:0] out_417;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_417 (
            .in(out_416),
            .outp(out_417)
        );
        

        logic [WIDTH-1:0] out_418;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_418 (
            .a(out_355),
            .b(out_417),
            .outp(out_418)
        );        
        

        logic [WIDTH-1:0] out_419;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_419 (
            .in(out_418),
            .outp(out_419)
        );
        

        logic [WIDTH-1:0] out_420;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_420 (
            .a(out_9),
            .b(out_419),
            .outp(out_420)
        );        
        

        logic [WIDTH-1:0] out_421;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_421 (
            .a(out_414),
            .b(out_420),
            .outp(out_421)
        );        
        

        logic [WIDTH-1:0] out_422;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_422 (
            .a(out_419),
            .b(out_21),
            .outp(out_422)
        );        
        

        logic [WIDTH-1:0] out_423;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_423 (
            .a(out_421),
            .b(out_422),
            .outp(out_423)
        );        
        

        logic [WIDTH-1:0] out_424;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_424 (
            .a(out_411),
            .b(out_423),
            .outp(out_424)
        );        
        

        logic [WIDTH-1:0] out_425;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6205)
        ) inst_425 (
            .outp(out_425)
        );
        

        logic [WIDTH-1:0] out_426;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_426 (
            .a(out_3),
            .b(out_425),
            .outp(out_426)
        );        
        

        logic [WIDTH-1:0] out_427;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_427 (
            .in(out_426),
            .outp(out_427)
        );
        

        logic [WIDTH-1:0] out_428;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_428 (
            .a(out_355),
            .b(out_427),
            .outp(out_428)
        );        
        

        logic [WIDTH-1:0] out_429;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_429 (
            .in(out_428),
            .outp(out_429)
        );
        

        logic [WIDTH-1:0] out_430;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_430 (
            .a(out_9),
            .b(out_429),
            .outp(out_430)
        );        
        

        logic [WIDTH-1:0] out_431;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_431 (
            .a(out_429),
            .b(out_21),
            .outp(out_431)
        );        
        

        logic [WIDTH-1:0] out_432;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_432 (
            .a(out_430),
            .b(out_431),
            .outp(out_432)
        );        
        

        logic [WIDTH-1:0] out_433;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_433 (
            .a(out_424),
            .b(out_432),
            .outp(out_433)
        );        
        

        logic [WIDTH-1:0] out_434;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.142001)
        ) inst_434 (
            .outp(out_434)
        );
        

        logic [WIDTH-1:0] out_435;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_435 (
            .a(out_434),
            .b(out_3),
            .outp(out_435)
        );        
        

        logic [WIDTH-1:0] out_436;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_436 (
            .a(out_94),
            .b(out_435),
            .outp(out_436)
        );        
        

        logic [WIDTH-1:0] out_437;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.242001)
        ) inst_437 (
            .outp(out_437)
        );
        

        logic [WIDTH-1:0] out_438;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_438 (
            .a(out_437),
            .b(out_3),
            .outp(out_438)
        );        
        

        logic [WIDTH-1:0] out_439;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_439 (
            .in(out_438),
            .outp(out_439)
        );
        

        logic [WIDTH-1:0] out_440;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_440 (
            .a(out_436),
            .b(out_439),
            .outp(out_440)
        );        
        

        logic [WIDTH-1:0] out_441;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.85)
        ) inst_441 (
            .outp(out_441)
        );
        

        logic [WIDTH-1:0] out_442;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_442 (
            .a(out_441),
            .b(out_14),
            .outp(out_442)
        );        
        

        logic [WIDTH-1:0] out_443;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_443 (
            .a(out_440),
            .b(out_442),
            .outp(out_443)
        );        
        

        logic [WIDTH-1:0] out_444;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_444 (
            .a(out_433),
            .b(out_443),
            .outp(out_444)
        );        
        

        logic [WIDTH-1:0] out_445;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.392001)
        ) inst_445 (
            .outp(out_445)
        );
        

        logic [WIDTH-1:0] out_446;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_446 (
            .a(out_445),
            .b(out_3),
            .outp(out_446)
        );        
        

        logic [WIDTH-1:0] out_447;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_447 (
            .a(out_94),
            .b(out_446),
            .outp(out_447)
        );        
        

        logic [WIDTH-1:0] out_448;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.492001)
        ) inst_448 (
            .outp(out_448)
        );
        

        logic [WIDTH-1:0] out_449;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_449 (
            .a(out_448),
            .b(out_3),
            .outp(out_449)
        );        
        

        logic [WIDTH-1:0] out_450;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_450 (
            .in(out_449),
            .outp(out_450)
        );
        

        logic [WIDTH-1:0] out_451;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_451 (
            .a(out_447),
            .b(out_450),
            .outp(out_451)
        );        
        

        logic [WIDTH-1:0] out_452;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.675)
        ) inst_452 (
            .outp(out_452)
        );
        

        logic [WIDTH-1:0] out_453;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_453 (
            .a(out_452),
            .b(out_14),
            .outp(out_453)
        );        
        

        logic [WIDTH-1:0] out_454;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_454 (
            .a(out_451),
            .b(out_453),
            .outp(out_454)
        );        
        

        logic [WIDTH-1:0] out_455;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_455 (
            .a(out_444),
            .b(out_454),
            .outp(out_455)
        );        
        

        logic [WIDTH-1:0] out_456;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_456 (
            .a(out_323),
            .b(out_450),
            .outp(out_456)
        );        
        

        logic [WIDTH-1:0] out_457;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.157999)
        ) inst_457 (
            .outp(out_457)
        );
        

        logic [WIDTH-1:0] out_458;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_458 (
            .a(out_3),
            .b(out_457),
            .outp(out_458)
        );        
        

        logic [WIDTH-1:0] out_459;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_459 (
            .a(out_456),
            .b(out_458),
            .outp(out_459)
        );        
        

        logic [WIDTH-1:0] out_460;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.075)
        ) inst_460 (
            .outp(out_460)
        );
        

        logic [WIDTH-1:0] out_461;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0670004)
        ) inst_461 (
            .outp(out_461)
        );
        

        logic [WIDTH-1:0] out_462;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_462 (
            .a(out_461),
            .b(out_3),
            .outp(out_462)
        );        
        

        logic [WIDTH-1:0] out_463;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_463 (
            .in(out_462),
            .outp(out_463)
        );
        

        logic [WIDTH-1:0] out_464;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_464 (
            .in(out_442),
            .outp(out_464)
        );
        

        logic [WIDTH-1:0] out_465;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_465 (
            .a(out_463),
            .b(out_464),
            .outp(out_465)
        );        
        

        logic [WIDTH-1:0] out_466;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_466 (
            .in(out_465),
            .outp(out_466)
        );
        

        logic [WIDTH-1:0] out_467;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_467 (
            .a(out_460),
            .b(out_466),
            .outp(out_467)
        );        
        

        logic [WIDTH-1:0] out_468;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_468 (
            .a(out_466),
            .b(out_9),
            .outp(out_468)
        );        
        

        logic [WIDTH-1:0] out_469;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_469 (
            .a(out_467),
            .b(out_468),
            .outp(out_469)
        );        
        

        logic [WIDTH-1:0] out_470;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.317)
        ) inst_470 (
            .outp(out_470)
        );
        

        logic [WIDTH-1:0] out_471;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_471 (
            .a(out_470),
            .b(out_3),
            .outp(out_471)
        );        
        

        logic [WIDTH-1:0] out_472;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_472 (
            .in(out_471),
            .outp(out_472)
        );
        

        logic [WIDTH-1:0] out_473;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_473 (
            .a(out_472),
            .b(out_464),
            .outp(out_473)
        );        
        

        logic [WIDTH-1:0] out_474;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_474 (
            .in(out_473),
            .outp(out_474)
        );
        

        logic [WIDTH-1:0] out_475;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_475 (
            .a(out_460),
            .b(out_474),
            .outp(out_475)
        );        
        

        logic [WIDTH-1:0] out_476;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_476 (
            .a(out_474),
            .b(out_9),
            .outp(out_476)
        );        
        

        logic [WIDTH-1:0] out_477;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_477 (
            .a(out_475),
            .b(out_476),
            .outp(out_477)
        );        
        

        logic [WIDTH-1:0] out_478;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_478 (
            .a(out_469),
            .b(out_477),
            .outp(out_478)
        );        
        

        logic [WIDTH-1:0] out_479;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_479 (
            .a(out_459),
            .b(out_478),
            .outp(out_479)
        );        
        

        logic [WIDTH-1:0] out_480;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.85)
        ) inst_480 (
            .outp(out_480)
        );
        

        logic [WIDTH-1:0] out_481;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_481 (
            .a(out_480),
            .b(out_14),
            .outp(out_481)
        );        
        

        logic [WIDTH-1:0] out_482;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_482 (
            .in(out_481),
            .outp(out_482)
        );
        

        logic [WIDTH-1:0] out_483;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_483 (
            .a(out_479),
            .b(out_482),
            .outp(out_483)
        );        
        

        logic [WIDTH-1:0] out_484;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_484 (
            .a(out_455),
            .b(out_483),
            .outp(out_484)
        );        
        

        logic [WIDTH-1:0] out_485;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.592)
        ) inst_485 (
            .outp(out_485)
        );
        

        logic [WIDTH-1:0] out_486;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_486 (
            .a(out_485),
            .b(out_3),
            .outp(out_486)
        );        
        

        logic [WIDTH-1:0] out_487;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_487 (
            .a(out_372),
            .b(out_486),
            .outp(out_487)
        );        
        

        logic [WIDTH-1:0] out_488;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.692001)
        ) inst_488 (
            .outp(out_488)
        );
        

        logic [WIDTH-1:0] out_489;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_489 (
            .a(out_488),
            .b(out_3),
            .outp(out_489)
        );        
        

        logic [WIDTH-1:0] out_490;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_490 (
            .in(out_489),
            .outp(out_490)
        );
        

        logic [WIDTH-1:0] out_491;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_491 (
            .a(out_487),
            .b(out_490),
            .outp(out_491)
        );        
        

        logic [WIDTH-1:0] out_492;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_492 (
            .a(out_484),
            .b(out_491),
            .outp(out_492)
        );        
        

        logic [WIDTH-1:0] out_493;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.042)
        ) inst_493 (
            .outp(out_493)
        );
        

        logic [WIDTH-1:0] out_494;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_494 (
            .a(out_493),
            .b(out_3),
            .outp(out_494)
        );        
        

        logic [WIDTH-1:0] out_495;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_495 (
            .a(out_404),
            .b(out_494),
            .outp(out_495)
        );        
        

        logic [WIDTH-1:0] out_496;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.142)
        ) inst_496 (
            .outp(out_496)
        );
        

        logic [WIDTH-1:0] out_497;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_497 (
            .a(out_496),
            .b(out_3),
            .outp(out_497)
        );        
        

        logic [WIDTH-1:0] out_498;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_498 (
            .in(out_497),
            .outp(out_498)
        );
        

        logic [WIDTH-1:0] out_499;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_499 (
            .a(out_495),
            .b(out_498),
            .outp(out_499)
        );        
        

        logic [WIDTH-1:0] out_500;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_500 (
            .a(out_492),
            .b(out_499),
            .outp(out_500)
        );        
        

        logic [WIDTH-1:0] out_501;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_501 (
            .a(out_412),
            .b(out_486),
            .outp(out_501)
        );        
        

        logic [WIDTH-1:0] out_502;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_502 (
            .a(out_501),
            .b(out_498),
            .outp(out_502)
        );        
        

        logic [WIDTH-1:0] out_503;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.867001)
        ) inst_503 (
            .outp(out_503)
        );
        

        logic [WIDTH-1:0] out_504;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_504 (
            .a(out_503),
            .b(out_3),
            .outp(out_504)
        );        
        

        logic [WIDTH-1:0] out_505;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_505 (
            .in(out_504),
            .outp(out_505)
        );
        

        logic [WIDTH-1:0] out_506;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_506 (
            .a(out_355),
            .b(out_505),
            .outp(out_506)
        );        
        

        logic [WIDTH-1:0] out_507;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_507 (
            .in(out_506),
            .outp(out_507)
        );
        

        logic [WIDTH-1:0] out_508;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_508 (
            .a(out_9),
            .b(out_507),
            .outp(out_508)
        );        
        

        logic [WIDTH-1:0] out_509;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_509 (
            .a(out_502),
            .b(out_508),
            .outp(out_509)
        );        
        

        logic [WIDTH-1:0] out_510;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_510 (
            .a(out_507),
            .b(out_21),
            .outp(out_510)
        );        
        

        logic [WIDTH-1:0] out_511;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_511 (
            .a(out_509),
            .b(out_510),
            .outp(out_511)
        );        
        

        logic [WIDTH-1:0] out_512;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_512 (
            .a(out_500),
            .b(out_511),
            .outp(out_512)
        );        
        

        logic [WIDTH-1:0] out_513;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.267)
        ) inst_513 (
            .outp(out_513)
        );
        

        logic [WIDTH-1:0] out_514;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_514 (
            .a(out_513),
            .b(out_3),
            .outp(out_514)
        );        
        

        logic [WIDTH-1:0] out_515;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_515 (
            .a(out_95),
            .b(out_514),
            .outp(out_515)
        );        
        

        logic [WIDTH-1:0] out_516;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.367)
        ) inst_516 (
            .outp(out_516)
        );
        

        logic [WIDTH-1:0] out_517;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_517 (
            .a(out_516),
            .b(out_3),
            .outp(out_517)
        );        
        

        logic [WIDTH-1:0] out_518;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_518 (
            .in(out_517),
            .outp(out_518)
        );
        

        logic [WIDTH-1:0] out_519;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_519 (
            .a(out_515),
            .b(out_518),
            .outp(out_519)
        );        
        

        logic [WIDTH-1:0] out_520;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_520 (
            .a(out_512),
            .b(out_519),
            .outp(out_520)
        );        
        

        logic [WIDTH-1:0] out_521;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.575)
        ) inst_521 (
            .outp(out_521)
        );
        

        logic [WIDTH-1:0] out_522;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_522 (
            .a(out_521),
            .b(out_14),
            .outp(out_522)
        );        
        

        logic [WIDTH-1:0] out_523;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_523 (
            .in(out_522),
            .outp(out_523)
        );
        

        logic [WIDTH-1:0] out_524;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_524 (
            .a(out_104),
            .b(out_523),
            .outp(out_524)
        );        
        

        logic [WIDTH-1:0] out_525;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.942)
        ) inst_525 (
            .outp(out_525)
        );
        

        logic [WIDTH-1:0] out_526;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_526 (
            .a(out_525),
            .b(out_3),
            .outp(out_526)
        );        
        

        logic [WIDTH-1:0] out_527;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_527 (
            .a(out_524),
            .b(out_526),
            .outp(out_527)
        );        
        

        logic [WIDTH-1:0] out_528;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.042)
        ) inst_528 (
            .outp(out_528)
        );
        

        logic [WIDTH-1:0] out_529;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_529 (
            .a(out_528),
            .b(out_3),
            .outp(out_529)
        );        
        

        logic [WIDTH-1:0] out_530;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_530 (
            .in(out_529),
            .outp(out_530)
        );
        

        logic [WIDTH-1:0] out_531;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_531 (
            .a(out_527),
            .b(out_530),
            .outp(out_531)
        );        
        

        logic [WIDTH-1:0] out_532;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_532 (
            .a(out_520),
            .b(out_531),
            .outp(out_532)
        );        
        

        logic [WIDTH-1:0] out_533;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.885)
        ) inst_533 (
            .outp(out_533)
        );
        

        logic [WIDTH-1:0] out_534;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_534 (
            .a(out_533),
            .b(out_14),
            .outp(out_534)
        );        
        

        logic [WIDTH-1:0] out_535;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.975)
        ) inst_535 (
            .outp(out_535)
        );
        

        logic [WIDTH-1:0] out_536;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_536 (
            .a(out_535),
            .b(out_14),
            .outp(out_536)
        );        
        

        logic [WIDTH-1:0] out_537;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_537 (
            .in(out_536),
            .outp(out_537)
        );
        

        logic [WIDTH-1:0] out_538;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_538 (
            .a(out_534),
            .b(out_537),
            .outp(out_538)
        );        
        

        logic [WIDTH-1:0] out_539;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.458)
        ) inst_539 (
            .outp(out_539)
        );
        

        logic [WIDTH-1:0] out_540;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_540 (
            .a(out_3),
            .b(out_539),
            .outp(out_540)
        );        
        

        logic [WIDTH-1:0] out_541;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_541 (
            .a(out_538),
            .b(out_540),
            .outp(out_541)
        );        
        

        logic [WIDTH-1:0] out_542;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.958001)
        ) inst_542 (
            .outp(out_542)
        );
        

        logic [WIDTH-1:0] out_543;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_543 (
            .a(out_542),
            .b(out_3),
            .outp(out_543)
        );        
        

        logic [WIDTH-1:0] out_544;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_544 (
            .a(out_541),
            .b(out_543),
            .outp(out_544)
        );        
        

        logic [WIDTH-1:0] out_545;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.183)
        ) inst_545 (
            .outp(out_545)
        );
        

        logic [WIDTH-1:0] out_546;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_546 (
            .a(out_3),
            .b(out_545),
            .outp(out_546)
        );        
        

        logic [WIDTH-1:0] out_547;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_547 (
            .in(out_546),
            .outp(out_547)
        );
        

        logic [WIDTH-1:0] out_548;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_548 (
            .a(out_355),
            .b(out_547),
            .outp(out_548)
        );        
        

        logic [WIDTH-1:0] out_549;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_549 (
            .in(out_548),
            .outp(out_549)
        );
        

        logic [WIDTH-1:0] out_550;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_550 (
            .a(out_549),
            .b(out_21),
            .outp(out_550)
        );        
        

        logic [WIDTH-1:0] out_551;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.20125)
        ) inst_551 (
            .outp(out_551)
        );
        

        logic [WIDTH-1:0] out_552;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.28455)
        ) inst_552 (
            .outp(out_552)
        );
        

        logic [WIDTH-1:0] out_553;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_553 (
            .a(out_13),
            .b(out_552),
            .outp(out_553)
        );        
        

        logic [WIDTH-1:0] out_554;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_554 (
            .a(out_551),
            .b(out_553),
            .outp(out_554)
        );        
        

        logic [WIDTH-1:0] out_555;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.23577)
        ) inst_555 (
            .outp(out_555)
        );
        

        logic [WIDTH-1:0] out_556;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_556 (
            .a(out_1),
            .b(out_555),
            .outp(out_556)
        );        
        

        logic [WIDTH-1:0] out_557;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.1947)
        ) inst_557 (
            .outp(out_557)
        );
        

        logic [WIDTH-1:0] out_558;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.21951)
        ) inst_558 (
            .outp(out_558)
        );
        

        logic [WIDTH-1:0] out_559;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_559 (
            .a(out_13),
            .b(out_558),
            .outp(out_559)
        );        
        

        logic [WIDTH-1:0] out_560;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_560 (
            .a(out_557),
            .b(out_559),
            .outp(out_560)
        );        
        

        logic [WIDTH-1:0] out_561;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_561 (
            .a(out_556),
            .b(out_560),
            .outp(out_561)
        );        
        

        logic [WIDTH-1:0] out_562;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_562 (
            .a(out_554),
            .b(out_561),
            .outp(out_562)
        );        
        

        logic [WIDTH-1:0] out_563;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.1853)
        ) inst_563 (
            .outp(out_563)
        );
        

        logic [WIDTH-1:0] out_564;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_564 (
            .a(out_563),
            .b(out_556),
            .outp(out_564)
        );        
        

        logic [WIDTH-1:0] out_565;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.06504)
        ) inst_565 (
            .outp(out_565)
        );
        

        logic [WIDTH-1:0] out_566;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_566 (
            .a(out_13),
            .b(out_565),
            .outp(out_566)
        );        
        

        logic [WIDTH-1:0] out_567;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_567 (
            .a(out_564),
            .b(out_566),
            .outp(out_567)
        );        
        

        logic [WIDTH-1:0] out_568;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_568 (
            .in(out_567),
            .outp(out_568)
        );
        

        logic [WIDTH-1:0] out_569;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_569 (
            .a(out_562),
            .b(out_568),
            .outp(out_569)
        );        
        

        logic [WIDTH-1:0] out_570;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.1853)
        ) inst_570 (
            .outp(out_570)
        );
        

        logic [WIDTH-1:0] out_571;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_571 (
            .a(out_570),
            .b(out_556),
            .outp(out_571)
        );        
        

        logic [WIDTH-1:0] out_572;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_572 (
            .a(out_571),
            .b(out_566),
            .outp(out_572)
        );        
        

        logic [WIDTH-1:0] out_573;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_573 (
            .a(out_560),
            .b(out_556),
            .outp(out_573)
        );        
        

        logic [WIDTH-1:0] out_574;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_574 (
            .a(out_572),
            .b(out_573),
            .outp(out_574)
        );        
        

        logic [WIDTH-1:0] out_575;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_575 (
            .in(out_554),
            .outp(out_575)
        );
        

        logic [WIDTH-1:0] out_576;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_576 (
            .a(out_574),
            .b(out_575),
            .outp(out_576)
        );        
        

        logic [WIDTH-1:0] out_577;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_577 (
            .a(out_569),
            .b(out_576),
            .outp(out_577)
        );        
        

        logic [WIDTH-1:0] out_578;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_578 (
            .in(out_577),
            .outp(out_578)
        );
        

        logic [WIDTH-1:0] out_579;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_579 (
            .a(out_550),
            .b(out_578),
            .outp(out_579)
        );        
        

        logic [WIDTH-1:0] out_580;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_580 (
            .a(out_9),
            .b(out_549),
            .outp(out_580)
        );        
        

        logic [WIDTH-1:0] out_581;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_581 (
            .a(out_579),
            .b(out_580),
            .outp(out_581)
        );        
        

        logic [WIDTH-1:0] out_582;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_582 (
            .a(out_544),
            .b(out_581),
            .outp(out_582)
        );        
        

        logic [WIDTH-1:0] out_583;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_583 (
            .a(out_550),
            .b(out_582),
            .outp(out_583)
        );        
        

        logic [WIDTH-1:0] out_584;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_584 (
            .a(out_532),
            .b(out_583),
            .outp(out_584)
        );        
        

        logic [WIDTH-1:0] out_585;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_585 (
            .a(out_94),
            .b(out_442),
            .outp(out_585)
        );        
        

        logic [WIDTH-1:0] out_586;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.808001)
        ) inst_586 (
            .outp(out_586)
        );
        

        logic [WIDTH-1:0] out_587;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_587 (
            .a(out_3),
            .b(out_586),
            .outp(out_587)
        );        
        

        logic [WIDTH-1:0] out_588;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_588 (
            .a(out_585),
            .b(out_587),
            .outp(out_588)
        );        
        

        logic [WIDTH-1:0] out_589;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.708)
        ) inst_589 (
            .outp(out_589)
        );
        

        logic [WIDTH-1:0] out_590;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_590 (
            .a(out_589),
            .b(out_3),
            .outp(out_590)
        );        
        

        logic [WIDTH-1:0] out_591;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_591 (
            .a(out_588),
            .b(out_590),
            .outp(out_591)
        );        
        

        logic [WIDTH-1:0] out_592;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_592 (
            .a(out_584),
            .b(out_591),
            .outp(out_592)
        );        
        

        logic [WIDTH-1:0] out_593;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.558001)
        ) inst_593 (
            .outp(out_593)
        );
        

        logic [WIDTH-1:0] out_594;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_594 (
            .a(out_3),
            .b(out_593),
            .outp(out_594)
        );        
        

        logic [WIDTH-1:0] out_595;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_595 (
            .a(out_585),
            .b(out_594),
            .outp(out_595)
        );        
        

        logic [WIDTH-1:0] out_596;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.458)
        ) inst_596 (
            .outp(out_596)
        );
        

        logic [WIDTH-1:0] out_597;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_597 (
            .a(out_596),
            .b(out_3),
            .outp(out_597)
        );        
        

        logic [WIDTH-1:0] out_598;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_598 (
            .a(out_595),
            .b(out_597),
            .outp(out_598)
        );        
        

        logic [WIDTH-1:0] out_599;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_599 (
            .a(out_592),
            .b(out_598),
            .outp(out_599)
        );        
        

        logic [WIDTH-1:0] out_600;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_600 (
            .a(out_94),
            .b(out_453),
            .outp(out_600)
        );        
        

        logic [WIDTH-1:0] out_601;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.308001)
        ) inst_601 (
            .outp(out_601)
        );
        

        logic [WIDTH-1:0] out_602;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_602 (
            .a(out_3),
            .b(out_601),
            .outp(out_602)
        );        
        

        logic [WIDTH-1:0] out_603;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_603 (
            .a(out_600),
            .b(out_602),
            .outp(out_603)
        );        
        

        logic [WIDTH-1:0] out_604;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.208)
        ) inst_604 (
            .outp(out_604)
        );
        

        logic [WIDTH-1:0] out_605;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_605 (
            .a(out_604),
            .b(out_3),
            .outp(out_605)
        );        
        

        logic [WIDTH-1:0] out_606;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_606 (
            .a(out_603),
            .b(out_605),
            .outp(out_606)
        );        
        

        logic [WIDTH-1:0] out_607;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_607 (
            .a(out_599),
            .b(out_606),
            .outp(out_607)
        );        
        

        logic [WIDTH-1:0] out_608;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_608 (
            .a(out_323),
            .b(out_605),
            .outp(out_608)
        );        
        

        logic [WIDTH-1:0] out_609;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_609 (
            .a(out_608),
            .b(out_482),
            .outp(out_609)
        );        
        

        logic [WIDTH-1:0] out_610;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.858)
        ) inst_610 (
            .outp(out_610)
        );
        

        logic [WIDTH-1:0] out_611;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_611 (
            .a(out_3),
            .b(out_610),
            .outp(out_611)
        );        
        

        logic [WIDTH-1:0] out_612;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_612 (
            .a(out_609),
            .b(out_611),
            .outp(out_612)
        );        
        

        logic [WIDTH-1:0] out_613;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.633)
        ) inst_613 (
            .outp(out_613)
        );
        

        logic [WIDTH-1:0] out_614;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_614 (
            .a(out_3),
            .b(out_613),
            .outp(out_614)
        );        
        

        logic [WIDTH-1:0] out_615;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_615 (
            .in(out_614),
            .outp(out_615)
        );
        

        logic [WIDTH-1:0] out_616;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_616 (
            .a(out_464),
            .b(out_615),
            .outp(out_616)
        );        
        

        logic [WIDTH-1:0] out_617;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_617 (
            .in(out_616),
            .outp(out_617)
        );
        

        logic [WIDTH-1:0] out_618;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_618 (
            .a(out_460),
            .b(out_617),
            .outp(out_618)
        );        
        

        logic [WIDTH-1:0] out_619;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_619 (
            .a(out_617),
            .b(out_9),
            .outp(out_619)
        );        
        

        logic [WIDTH-1:0] out_620;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_620 (
            .a(out_618),
            .b(out_619),
            .outp(out_620)
        );        
        

        logic [WIDTH-1:0] out_621;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.383)
        ) inst_621 (
            .outp(out_621)
        );
        

        logic [WIDTH-1:0] out_622;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_622 (
            .a(out_3),
            .b(out_621),
            .outp(out_622)
        );        
        

        logic [WIDTH-1:0] out_623;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_623 (
            .in(out_622),
            .outp(out_623)
        );
        

        logic [WIDTH-1:0] out_624;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_624 (
            .a(out_464),
            .b(out_623),
            .outp(out_624)
        );        
        

        logic [WIDTH-1:0] out_625;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_625 (
            .in(out_624),
            .outp(out_625)
        );
        

        logic [WIDTH-1:0] out_626;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_626 (
            .a(out_460),
            .b(out_625),
            .outp(out_626)
        );        
        

        logic [WIDTH-1:0] out_627;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_627 (
            .a(out_625),
            .b(out_9),
            .outp(out_627)
        );        
        

        logic [WIDTH-1:0] out_628;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_628 (
            .a(out_626),
            .b(out_627),
            .outp(out_628)
        );        
        

        logic [WIDTH-1:0] out_629;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_629 (
            .a(out_620),
            .b(out_628),
            .outp(out_629)
        );        
        

        logic [WIDTH-1:0] out_630;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_630 (
            .a(out_612),
            .b(out_629),
            .outp(out_630)
        );        
        

        logic [WIDTH-1:0] out_631;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_631 (
            .a(out_607),
            .b(out_630),
            .outp(out_631)
        );        
        

        logic [WIDTH-1:0] out_632;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.108)
        ) inst_632 (
            .outp(out_632)
        );
        

        logic [WIDTH-1:0] out_633;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_633 (
            .a(out_3),
            .b(out_632),
            .outp(out_633)
        );        
        

        logic [WIDTH-1:0] out_634;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_634 (
            .a(out_585),
            .b(out_633),
            .outp(out_634)
        );        
        

        logic [WIDTH-1:0] out_635;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.00799942)
        ) inst_635 (
            .outp(out_635)
        );
        

        logic [WIDTH-1:0] out_636;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_636 (
            .a(out_635),
            .b(out_3),
            .outp(out_636)
        );        
        

        logic [WIDTH-1:0] out_637;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_637 (
            .a(out_634),
            .b(out_636),
            .outp(out_637)
        );        
        

        logic [WIDTH-1:0] out_638;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_638 (
            .a(out_631),
            .b(out_637),
            .outp(out_638)
        );        
        

        logic [WIDTH-1:0] out_639;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.767)
        ) inst_639 (
            .outp(out_639)
        );
        

        logic [WIDTH-1:0] out_640;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_640 (
            .a(out_639),
            .b(out_3),
            .outp(out_640)
        );        
        

        logic [WIDTH-1:0] out_641;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_641 (
            .in(out_640),
            .outp(out_641)
        );
        

        logic [WIDTH-1:0] out_642;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_642 (
            .a(out_355),
            .b(out_641),
            .outp(out_642)
        );        
        

        logic [WIDTH-1:0] out_643;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_643 (
            .in(out_642),
            .outp(out_643)
        );
        

        logic [WIDTH-1:0] out_644;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_644 (
            .a(out_9),
            .b(out_643),
            .outp(out_644)
        );        
        

        logic [WIDTH-1:0] out_645;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_645 (
            .a(out_643),
            .b(out_21),
            .outp(out_645)
        );        
        

        logic [WIDTH-1:0] out_646;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_646 (
            .a(out_644),
            .b(out_645),
            .outp(out_646)
        );        
        

        logic [WIDTH-1:0] out_647;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_647 (
            .a(out_638),
            .b(out_646),
            .outp(out_647)
        );        
        

        logic [WIDTH-1:0] out_648;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.13)
        ) inst_648 (
            .outp(out_648)
        );
        

        logic [WIDTH-1:0] out_649;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_649 (
            .a(out_124),
            .b(out_648),
            .outp(out_649)
        );        
        

        logic [WIDTH-1:0] out_650;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_650 (
            .a(out_649),
            .b(out_127),
            .outp(out_650)
        );        
        

        logic [WIDTH-1:0] out_651;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.52)
        ) inst_651 (
            .outp(out_651)
        );
        

        logic [WIDTH-1:0] out_652;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_652 (
            .a(out_651),
            .b(out_152),
            .outp(out_652)
        );        
        

        logic [WIDTH-1:0] out_653;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_653 (
            .in(out_652),
            .outp(out_653)
        );
        

        logic [WIDTH-1:0] out_654;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_654 (
            .a(out_650),
            .b(out_653),
            .outp(out_654)
        );        
        

        logic [WIDTH-1:0] out_655;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.665)
        ) inst_655 (
            .outp(out_655)
        );
        

        logic [WIDTH-1:0] out_656;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_656 (
            .a(out_131),
            .b(out_655),
            .outp(out_656)
        );        
        

        logic [WIDTH-1:0] out_657;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_657 (
            .a(out_656),
            .b(out_127),
            .outp(out_657)
        );        
        

        logic [WIDTH-1:0] out_658;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_658 (
            .in(out_657),
            .outp(out_658)
        );
        

        logic [WIDTH-1:0] out_659;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_659 (
            .a(out_654),
            .b(out_658),
            .outp(out_659)
        );        
        

        logic [WIDTH-1:0] out_660;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_660 (
            .a(out_647),
            .b(out_659),
            .outp(out_660)
        );        
        

        logic [WIDTH-1:0] out_661;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_661 (
            .in(out_650),
            .outp(out_661)
        );
        

        logic [WIDTH-1:0] out_662;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_662 (
            .a(out_661),
            .b(out_652),
            .outp(out_662)
        );        
        

        logic [WIDTH-1:0] out_663;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_663 (
            .a(out_662),
            .b(out_657),
            .outp(out_663)
        );        
        

        logic [WIDTH-1:0] out_664;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_664 (
            .a(out_660),
            .b(out_663),
            .outp(out_664)
        );        
        

        logic [WIDTH-1:0] out_665;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.61)
        ) inst_665 (
            .outp(out_665)
        );
        

        logic [WIDTH-1:0] out_666;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_666 (
            .a(out_131),
            .b(out_665),
            .outp(out_666)
        );        
        

        logic [WIDTH-1:0] out_667;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_667 (
            .a(out_666),
            .b(out_127),
            .outp(out_667)
        );        
        

        logic [WIDTH-1:0] out_668;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_668 (
            .a(out_661),
            .b(out_667),
            .outp(out_668)
        );        
        

        logic [WIDTH-1:0] out_669;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.465)
        ) inst_669 (
            .outp(out_669)
        );
        

        logic [WIDTH-1:0] out_670;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_670 (
            .a(out_669),
            .b(out_137),
            .outp(out_670)
        );        
        

        logic [WIDTH-1:0] out_671;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_671 (
            .a(out_668),
            .b(out_670),
            .outp(out_671)
        );        
        

        logic [WIDTH-1:0] out_672;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_672 (
            .a(out_664),
            .b(out_671),
            .outp(out_672)
        );        
        

        logic [WIDTH-1:0] out_673;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_673 (
            .in(out_667),
            .outp(out_673)
        );
        

        logic [WIDTH-1:0] out_674;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_674 (
            .a(out_650),
            .b(out_673),
            .outp(out_674)
        );        
        

        logic [WIDTH-1:0] out_675;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_675 (
            .in(out_670),
            .outp(out_675)
        );
        

        logic [WIDTH-1:0] out_676;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_676 (
            .a(out_674),
            .b(out_675),
            .outp(out_676)
        );        
        

        logic [WIDTH-1:0] out_677;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_677 (
            .a(out_672),
            .b(out_676),
            .outp(out_677)
        );        
        

        logic [WIDTH-1:0] out_678;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_678 (
            .a(out_103),
            .b(out_3),
            .outp(out_678)
        );        
        

        logic [WIDTH-1:0] out_679;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_679 (
            .a(out_538),
            .b(out_678),
            .outp(out_679)
        );        
        

        logic [WIDTH-1:0] out_680;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.15)
        ) inst_680 (
            .outp(out_680)
        );
        

        logic [WIDTH-1:0] out_681;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_681 (
            .a(out_680),
            .b(out_3),
            .outp(out_681)
        );        
        

        logic [WIDTH-1:0] out_682;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_682 (
            .in(out_681),
            .outp(out_682)
        );
        

        logic [WIDTH-1:0] out_683;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_683 (
            .a(out_679),
            .b(out_682),
            .outp(out_683)
        );        
        

        logic [WIDTH-1:0] out_684;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.925)
        ) inst_684 (
            .outp(out_684)
        );
        

        logic [WIDTH-1:0] out_685;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_685 (
            .a(out_684),
            .b(out_3),
            .outp(out_685)
        );        
        

        logic [WIDTH-1:0] out_686;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_686 (
            .in(out_685),
            .outp(out_686)
        );
        

        logic [WIDTH-1:0] out_687;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_687 (
            .a(out_355),
            .b(out_686),
            .outp(out_687)
        );        
        

        logic [WIDTH-1:0] out_688;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_688 (
            .in(out_687),
            .outp(out_688)
        );
        

        logic [WIDTH-1:0] out_689;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_689 (
            .a(out_688),
            .b(out_21),
            .outp(out_689)
        );        
        

        logic [WIDTH-1:0] out_690;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.485)
        ) inst_690 (
            .outp(out_690)
        );
        

        logic [WIDTH-1:0] out_691;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_691 (
            .a(out_690),
            .b(out_556),
            .outp(out_691)
        );        
        

        logic [WIDTH-1:0] out_692;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_692 (
            .a(out_691),
            .b(out_559),
            .outp(out_692)
        );        
        

        logic [WIDTH-1:0] out_693;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_693 (
            .a(out_554),
            .b(out_692),
            .outp(out_693)
        );        
        

        logic [WIDTH-1:0] out_694;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.865)
        ) inst_694 (
            .outp(out_694)
        );
        

        logic [WIDTH-1:0] out_695;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_695 (
            .a(out_556),
            .b(out_694),
            .outp(out_695)
        );        
        

        logic [WIDTH-1:0] out_696;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_696 (
            .a(out_695),
            .b(out_566),
            .outp(out_696)
        );        
        

        logic [WIDTH-1:0] out_697;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_697 (
            .in(out_696),
            .outp(out_697)
        );
        

        logic [WIDTH-1:0] out_698;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_698 (
            .a(out_693),
            .b(out_697),
            .outp(out_698)
        );        
        

        logic [WIDTH-1:0] out_699;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.865)
        ) inst_699 (
            .outp(out_699)
        );
        

        logic [WIDTH-1:0] out_700;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_700 (
            .a(out_556),
            .b(out_699),
            .outp(out_700)
        );        
        

        logic [WIDTH-1:0] out_701;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_701 (
            .a(out_700),
            .b(out_566),
            .outp(out_701)
        );        
        

        logic [WIDTH-1:0] out_702;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_702 (
            .a(out_575),
            .b(out_701),
            .outp(out_702)
        );        
        

        logic [WIDTH-1:0] out_703;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_703 (
            .a(out_559),
            .b(out_691),
            .outp(out_703)
        );        
        

        logic [WIDTH-1:0] out_704;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_704 (
            .a(out_702),
            .b(out_703),
            .outp(out_704)
        );        
        

        logic [WIDTH-1:0] out_705;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_705 (
            .a(out_698),
            .b(out_704),
            .outp(out_705)
        );        
        

        logic [WIDTH-1:0] out_706;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_706 (
            .in(out_705),
            .outp(out_706)
        );
        

        logic [WIDTH-1:0] out_707;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_707 (
            .a(out_689),
            .b(out_706),
            .outp(out_707)
        );        
        

        logic [WIDTH-1:0] out_708;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_708 (
            .a(out_9),
            .b(out_688),
            .outp(out_708)
        );        
        

        logic [WIDTH-1:0] out_709;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_709 (
            .a(out_707),
            .b(out_708),
            .outp(out_709)
        );        
        

        logic [WIDTH-1:0] out_710;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_710 (
            .a(out_683),
            .b(out_709),
            .outp(out_710)
        );        
        

        logic [WIDTH-1:0] out_711;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_711 (
            .a(out_689),
            .b(out_710),
            .outp(out_711)
        );        
        

        logic [WIDTH-1:0] out_712;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_712 (
            .a(out_677),
            .b(out_711),
            .outp(out_712)
        );        
        

        logic [WIDTH-1:0] out_713;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1)
        ) inst_713 (
            .outp(out_713)
        );
        

        logic [WIDTH-1:0] out_714;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_714 (
            .a(out_713),
            .b(out_14),
            .outp(out_714)
        );        
        

        logic [WIDTH-1:0] out_715;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.1)
        ) inst_715 (
            .outp(out_715)
        );
        

        logic [WIDTH-1:0] out_716;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_716 (
            .a(out_715),
            .b(out_14),
            .outp(out_716)
        );        
        

        logic [WIDTH-1:0] out_717;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_717 (
            .in(out_716),
            .outp(out_717)
        );
        

        logic [WIDTH-1:0] out_718;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_718 (
            .a(out_714),
            .b(out_717),
            .outp(out_718)
        );        
        

        logic [WIDTH-1:0] out_719;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.531)
        ) inst_719 (
            .outp(out_719)
        );
        

        logic [WIDTH-1:0] out_720;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_720 (
            .a(out_719),
            .b(out_3),
            .outp(out_720)
        );        
        

        logic [WIDTH-1:0] out_721;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_721 (
            .a(out_718),
            .b(out_720),
            .outp(out_721)
        );        
        

        logic [WIDTH-1:0] out_722;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.631)
        ) inst_722 (
            .outp(out_722)
        );
        

        logic [WIDTH-1:0] out_723;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_723 (
            .a(out_3),
            .b(out_722),
            .outp(out_723)
        );        
        

        logic [WIDTH-1:0] out_724;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_724 (
            .a(out_721),
            .b(out_723),
            .outp(out_724)
        );        
        

        logic [WIDTH-1:0] out_725;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_725 (
            .a(out_712),
            .b(out_724),
            .outp(out_725)
        );        
        

        logic [WIDTH-1:0] out_726;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.55)
        ) inst_726 (
            .outp(out_726)
        );
        

        logic [WIDTH-1:0] out_727;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_727 (
            .a(out_726),
            .b(out_14),
            .outp(out_727)
        );        
        

        logic [WIDTH-1:0] out_728;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.65)
        ) inst_728 (
            .outp(out_728)
        );
        

        logic [WIDTH-1:0] out_729;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_729 (
            .a(out_728),
            .b(out_14),
            .outp(out_729)
        );        
        

        logic [WIDTH-1:0] out_730;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_730 (
            .in(out_729),
            .outp(out_730)
        );
        

        logic [WIDTH-1:0] out_731;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_731 (
            .a(out_727),
            .b(out_730),
            .outp(out_731)
        );        
        

        logic [WIDTH-1:0] out_732;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.35601)
        ) inst_732 (
            .outp(out_732)
        );
        

        logic [WIDTH-1:0] out_733;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_733 (
            .a(out_732),
            .b(out_3),
            .outp(out_733)
        );        
        

        logic [WIDTH-1:0] out_734;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_734 (
            .a(out_731),
            .b(out_733),
            .outp(out_734)
        );        
        

        logic [WIDTH-1:0] out_735;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.531)
        ) inst_735 (
            .outp(out_735)
        );
        

        logic [WIDTH-1:0] out_736;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_736 (
            .a(out_3),
            .b(out_735),
            .outp(out_736)
        );        
        

        logic [WIDTH-1:0] out_737;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_737 (
            .a(out_734),
            .b(out_736),
            .outp(out_737)
        );        
        

        logic [WIDTH-1:0] out_738;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_738 (
            .a(out_725),
            .b(out_737),
            .outp(out_738)
        );        
        

        logic [WIDTH-1:0] out_739;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_739 (
            .a(out_717),
            .b(out_733),
            .outp(out_739)
        );        
        

        logic [WIDTH-1:0] out_740;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_740 (
            .a(out_739),
            .b(out_736),
            .outp(out_740)
        );        
        

        logic [WIDTH-1:0] out_741;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.0)
        ) inst_741 (
            .outp(out_741)
        );
        

        logic [WIDTH-1:0] out_742;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_742 (
            .a(out_741),
            .b(out_14),
            .outp(out_742)
        );        
        

        logic [WIDTH-1:0] out_743;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_743 (
            .a(out_740),
            .b(out_742),
            .outp(out_743)
        );        
        

        logic [WIDTH-1:0] out_744;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_744 (
            .a(out_738),
            .b(out_743),
            .outp(out_744)
        );        
        

        logic [WIDTH-1:0] out_745;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.631)
        ) inst_745 (
            .outp(out_745)
        );
        

        logic [WIDTH-1:0] out_746;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_746 (
            .a(out_745),
            .b(out_3),
            .outp(out_746)
        );        
        

        logic [WIDTH-1:0] out_747;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_747 (
            .a(out_718),
            .b(out_746),
            .outp(out_747)
        );        
        

        logic [WIDTH-1:0] out_748;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.356)
        ) inst_748 (
            .outp(out_748)
        );
        

        logic [WIDTH-1:0] out_749;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_749 (
            .a(out_3),
            .b(out_748),
            .outp(out_749)
        );        
        

        logic [WIDTH-1:0] out_750;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_750 (
            .a(out_747),
            .b(out_749),
            .outp(out_750)
        );        
        

        logic [WIDTH-1:0] out_751;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.825)
        ) inst_751 (
            .outp(out_751)
        );
        

        logic [WIDTH-1:0] out_752;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_752 (
            .a(out_751),
            .b(out_14),
            .outp(out_752)
        );        
        

        logic [WIDTH-1:0] out_753;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_753 (
            .in(out_752),
            .outp(out_753)
        );
        

        logic [WIDTH-1:0] out_754;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_754 (
            .in(out_733),
            .outp(out_754)
        );
        

        logic [WIDTH-1:0] out_755;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_755 (
            .a(out_753),
            .b(out_754),
            .outp(out_755)
        );        
        

        logic [WIDTH-1:0] out_756;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_756 (
            .in(out_755),
            .outp(out_756)
        );
        

        logic [WIDTH-1:0] out_757;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_757 (
            .a(out_9),
            .b(out_756),
            .outp(out_757)
        );        
        

        logic [WIDTH-1:0] out_758;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_758 (
            .a(out_750),
            .b(out_757),
            .outp(out_758)
        );        
        

        logic [WIDTH-1:0] out_759;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_759 (
            .a(out_756),
            .b(out_21),
            .outp(out_759)
        );        
        

        logic [WIDTH-1:0] out_760;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_760 (
            .a(out_758),
            .b(out_759),
            .outp(out_760)
        );        
        

        logic [WIDTH-1:0] out_761;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_761 (
            .a(out_744),
            .b(out_760),
            .outp(out_761)
        );        
        

        logic [WIDTH-1:0] out_762;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_762 (
            .a(out_713),
            .b(out_3),
            .outp(out_762)
        );        
        

        logic [WIDTH-1:0] out_763;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_763 (
            .a(out_372),
            .b(out_762),
            .outp(out_763)
        );        
        

        logic [WIDTH-1:0] out_764;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2)
        ) inst_764 (
            .outp(out_764)
        );
        

        logic [WIDTH-1:0] out_765;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_765 (
            .a(out_764),
            .b(out_3),
            .outp(out_765)
        );        
        

        logic [WIDTH-1:0] out_766;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_766 (
            .in(out_765),
            .outp(out_766)
        );
        

        logic [WIDTH-1:0] out_767;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_767 (
            .a(out_763),
            .b(out_766),
            .outp(out_767)
        );        
        

        logic [WIDTH-1:0] out_768;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_768 (
            .a(out_761),
            .b(out_767),
            .outp(out_768)
        );        
        

        logic [WIDTH-1:0] out_769;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.02143)
        ) inst_769 (
            .outp(out_769)
        );
        

        logic [WIDTH-1:0] out_770;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_770 (
            .a(out_769),
            .b(out_194),
            .outp(out_770)
        );        
        

        logic [WIDTH-1:0] out_771;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_771 (
            .a(out_372),
            .b(out_770),
            .outp(out_771)
        );        
        

        logic [WIDTH-1:0] out_772;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.57143)
        ) inst_772 (
            .outp(out_772)
        );
        

        logic [WIDTH-1:0] out_773;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_773 (
            .a(out_772),
            .b(out_194),
            .outp(out_773)
        );        
        

        logic [WIDTH-1:0] out_774;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_774 (
            .in(out_773),
            .outp(out_774)
        );
        

        logic [WIDTH-1:0] out_775;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_775 (
            .a(out_771),
            .b(out_774),
            .outp(out_775)
        );        
        

        logic [WIDTH-1:0] out_776;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_776 (
            .in(out_93),
            .outp(out_776)
        );
        

        logic [WIDTH-1:0] out_777;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.02679)
        ) inst_777 (
            .outp(out_777)
        );
        

        logic [WIDTH-1:0] out_778;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_778 (
            .a(out_777),
            .b(out_204),
            .outp(out_778)
        );        
        

        logic [WIDTH-1:0] out_779;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_779 (
            .in(out_778),
            .outp(out_779)
        );
        

        logic [WIDTH-1:0] out_780;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_780 (
            .a(out_776),
            .b(out_779),
            .outp(out_780)
        );        
        

        logic [WIDTH-1:0] out_781;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_781 (
            .in(out_780),
            .outp(out_781)
        );
        

        logic [WIDTH-1:0] out_782;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_782 (
            .a(out_200),
            .b(out_781),
            .outp(out_782)
        );        
        

        logic [WIDTH-1:0] out_783;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_783 (
            .a(out_775),
            .b(out_782),
            .outp(out_783)
        );        
        

        logic [WIDTH-1:0] out_784;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_784 (
            .in(out_770),
            .outp(out_784)
        );
        

        logic [WIDTH-1:0] out_785;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_785 (
            .a(out_776),
            .b(out_784),
            .outp(out_785)
        );        
        

        logic [WIDTH-1:0] out_786;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_786 (
            .in(out_785),
            .outp(out_786)
        );
        

        logic [WIDTH-1:0] out_787;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_787 (
            .a(out_786),
            .b(out_214),
            .outp(out_787)
        );        
        

        logic [WIDTH-1:0] out_788;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_788 (
            .a(out_783),
            .b(out_787),
            .outp(out_788)
        );        
        

        logic [WIDTH-1:0] out_789;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_789 (
            .a(out_768),
            .b(out_788),
            .outp(out_789)
        );        
        

        logic [WIDTH-1:0] out_790;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.3)
        ) inst_790 (
            .outp(out_790)
        );
        

        logic [WIDTH-1:0] out_791;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_791 (
            .a(out_790),
            .b(out_3),
            .outp(out_791)
        );        
        

        logic [WIDTH-1:0] out_792;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_792 (
            .a(out_538),
            .b(out_791),
            .outp(out_792)
        );        
        

        logic [WIDTH-1:0] out_793;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.8)
        ) inst_793 (
            .outp(out_793)
        );
        

        logic [WIDTH-1:0] out_794;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_794 (
            .a(out_793),
            .b(out_3),
            .outp(out_794)
        );        
        

        logic [WIDTH-1:0] out_795;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_795 (
            .in(out_794),
            .outp(out_795)
        );
        

        logic [WIDTH-1:0] out_796;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_796 (
            .a(out_792),
            .b(out_795),
            .outp(out_796)
        );        
        

        logic [WIDTH-1:0] out_797;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.575)
        ) inst_797 (
            .outp(out_797)
        );
        

        logic [WIDTH-1:0] out_798;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_798 (
            .a(out_797),
            .b(out_3),
            .outp(out_798)
        );        
        

        logic [WIDTH-1:0] out_799;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_799 (
            .in(out_798),
            .outp(out_799)
        );
        

        logic [WIDTH-1:0] out_800;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_800 (
            .a(out_355),
            .b(out_799),
            .outp(out_800)
        );        
        

        logic [WIDTH-1:0] out_801;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_801 (
            .in(out_800),
            .outp(out_801)
        );
        

        logic [WIDTH-1:0] out_802;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_802 (
            .a(out_801),
            .b(out_21),
            .outp(out_802)
        );        
        

        logic [WIDTH-1:0] out_803;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.11375)
        ) inst_803 (
            .outp(out_803)
        );
        

        logic [WIDTH-1:0] out_804;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_804 (
            .a(out_803),
            .b(out_556),
            .outp(out_804)
        );        
        

        logic [WIDTH-1:0] out_805;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_805 (
            .a(out_804),
            .b(out_559),
            .outp(out_805)
        );        
        

        logic [WIDTH-1:0] out_806;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_806 (
            .a(out_554),
            .b(out_805),
            .outp(out_806)
        );        
        

        logic [WIDTH-1:0] out_807;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.49375)
        ) inst_807 (
            .outp(out_807)
        );
        

        logic [WIDTH-1:0] out_808;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_808 (
            .a(out_556),
            .b(out_807),
            .outp(out_808)
        );        
        

        logic [WIDTH-1:0] out_809;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_809 (
            .a(out_808),
            .b(out_566),
            .outp(out_809)
        );        
        

        logic [WIDTH-1:0] out_810;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_810 (
            .in(out_809),
            .outp(out_810)
        );
        

        logic [WIDTH-1:0] out_811;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_811 (
            .a(out_806),
            .b(out_810),
            .outp(out_811)
        );        
        

        logic [WIDTH-1:0] out_812;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.49375)
        ) inst_812 (
            .outp(out_812)
        );
        

        logic [WIDTH-1:0] out_813;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_813 (
            .a(out_556),
            .b(out_812),
            .outp(out_813)
        );        
        

        logic [WIDTH-1:0] out_814;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_814 (
            .a(out_813),
            .b(out_566),
            .outp(out_814)
        );        
        

        logic [WIDTH-1:0] out_815;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_815 (
            .a(out_575),
            .b(out_814),
            .outp(out_815)
        );        
        

        logic [WIDTH-1:0] out_816;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_816 (
            .a(out_559),
            .b(out_804),
            .outp(out_816)
        );        
        

        logic [WIDTH-1:0] out_817;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_817 (
            .a(out_815),
            .b(out_816),
            .outp(out_817)
        );        
        

        logic [WIDTH-1:0] out_818;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_818 (
            .a(out_811),
            .b(out_817),
            .outp(out_818)
        );        
        

        logic [WIDTH-1:0] out_819;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_819 (
            .in(out_818),
            .outp(out_819)
        );
        

        logic [WIDTH-1:0] out_820;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_820 (
            .a(out_802),
            .b(out_819),
            .outp(out_820)
        );        
        

        logic [WIDTH-1:0] out_821;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_821 (
            .a(out_9),
            .b(out_801),
            .outp(out_821)
        );        
        

        logic [WIDTH-1:0] out_822;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_822 (
            .a(out_820),
            .b(out_821),
            .outp(out_822)
        );        
        

        logic [WIDTH-1:0] out_823;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_823 (
            .a(out_796),
            .b(out_822),
            .outp(out_823)
        );        
        

        logic [WIDTH-1:0] out_824;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_824 (
            .a(out_802),
            .b(out_823),
            .outp(out_824)
        );        
        

        logic [WIDTH-1:0] out_825;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_825 (
            .a(out_789),
            .b(out_824),
            .outp(out_825)
        );        
        

        logic [WIDTH-1:0] out_826;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.01)
        ) inst_826 (
            .outp(out_826)
        );
        

        logic [WIDTH-1:0] out_827;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_827 (
            .a(out_826),
            .b(out_127),
            .outp(out_827)
        );        
        

        logic [WIDTH-1:0] out_828;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_828 (
            .a(out_827),
            .b(out_131),
            .outp(out_828)
        );        
        

        logic [WIDTH-1:0] out_829;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_829 (
            .a(out_653),
            .b(out_828),
            .outp(out_829)
        );        
        

        logic [WIDTH-1:0] out_830;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.545)
        ) inst_830 (
            .outp(out_830)
        );
        

        logic [WIDTH-1:0] out_831;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_831 (
            .a(out_830),
            .b(out_127),
            .outp(out_831)
        );        
        

        logic [WIDTH-1:0] out_832;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_832 (
            .a(out_124),
            .b(out_831),
            .outp(out_832)
        );        
        

        logic [WIDTH-1:0] out_833;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_833 (
            .a(out_829),
            .b(out_832),
            .outp(out_833)
        );        
        

        logic [WIDTH-1:0] out_834;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_834 (
            .a(out_825),
            .b(out_833),
            .outp(out_834)
        );        
        

        logic [WIDTH-1:0] out_835;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_835 (
            .a(out_831),
            .b(out_124),
            .outp(out_835)
        );        
        

        logic [WIDTH-1:0] out_836;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_836 (
            .a(out_652),
            .b(out_835),
            .outp(out_836)
        );        
        

        logic [WIDTH-1:0] out_837;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_837 (
            .a(out_131),
            .b(out_827),
            .outp(out_837)
        );        
        

        logic [WIDTH-1:0] out_838;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_838 (
            .a(out_836),
            .b(out_837),
            .outp(out_838)
        );        
        

        logic [WIDTH-1:0] out_839;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_839 (
            .a(out_834),
            .b(out_838),
            .outp(out_839)
        );        
        

        logic [WIDTH-1:0] out_840;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_840 (
            .a(out_835),
            .b(out_670),
            .outp(out_840)
        );        
        

        logic [WIDTH-1:0] out_841;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.065)
        ) inst_841 (
            .outp(out_841)
        );
        

        logic [WIDTH-1:0] out_842;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_842 (
            .a(out_841),
            .b(out_127),
            .outp(out_842)
        );        
        

        logic [WIDTH-1:0] out_843;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_843 (
            .a(out_131),
            .b(out_842),
            .outp(out_843)
        );        
        

        logic [WIDTH-1:0] out_844;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_844 (
            .a(out_840),
            .b(out_843),
            .outp(out_844)
        );        
        

        logic [WIDTH-1:0] out_845;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_845 (
            .a(out_839),
            .b(out_844),
            .outp(out_845)
        );        
        

        logic [WIDTH-1:0] out_846;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_846 (
            .a(out_842),
            .b(out_131),
            .outp(out_846)
        );        
        

        logic [WIDTH-1:0] out_847;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_847 (
            .a(out_832),
            .b(out_846),
            .outp(out_847)
        );        
        

        logic [WIDTH-1:0] out_848;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_848 (
            .a(out_847),
            .b(out_675),
            .outp(out_848)
        );        
        

        logic [WIDTH-1:0] out_849;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_849 (
            .a(out_845),
            .b(out_848),
            .outp(out_849)
        );        
        

        logic [WIDTH-1:0] out_850;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.225)
        ) inst_850 (
            .outp(out_850)
        );
        

        logic [WIDTH-1:0] out_851;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_851 (
            .a(out_850),
            .b(out_14),
            .outp(out_851)
        );        
        

        logic [WIDTH-1:0] out_852;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_852 (
            .in(out_851),
            .outp(out_852)
        );
        

        logic [WIDTH-1:0] out_853;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.733)
        ) inst_853 (
            .outp(out_853)
        );
        

        logic [WIDTH-1:0] out_854;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_854 (
            .a(out_3),
            .b(out_853),
            .outp(out_854)
        );        
        

        logic [WIDTH-1:0] out_855;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_855 (
            .in(out_854),
            .outp(out_855)
        );
        

        logic [WIDTH-1:0] out_856;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_856 (
            .a(out_852),
            .b(out_855),
            .outp(out_856)
        );        
        

        logic [WIDTH-1:0] out_857;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_857 (
            .in(out_856),
            .outp(out_857)
        );
        

        logic [WIDTH-1:0] out_858;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_858 (
            .a(out_857),
            .b(out_460),
            .outp(out_858)
        );        
        

        logic [WIDTH-1:0] out_859;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_859 (
            .a(out_849),
            .b(out_858),
            .outp(out_859)
        );        
        

        logic [WIDTH-1:0] out_860;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.65)
        ) inst_860 (
            .outp(out_860)
        );
        

        logic [WIDTH-1:0] out_861;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_861 (
            .a(out_860),
            .b(out_566),
            .outp(out_861)
        );        
        

        logic [WIDTH-1:0] out_862;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_862 (
            .a(out_1),
            .b(out_565),
            .outp(out_862)
        );        
        

        logic [WIDTH-1:0] out_863;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.829)
        ) inst_863 (
            .outp(out_863)
        );
        

        logic [WIDTH-1:0] out_864;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_864 (
            .a(out_862),
            .b(out_863),
            .outp(out_864)
        );        
        

        logic [WIDTH-1:0] out_865;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_865 (
            .a(out_861),
            .b(out_864),
            .outp(out_865)
        );        
        

        logic [WIDTH-1:0] out_866;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0709989)
        ) inst_866 (
            .outp(out_866)
        );
        

        logic [WIDTH-1:0] out_867;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_867 (
            .a(out_1),
            .b(out_13),
            .outp(out_867)
        );        
        

        logic [WIDTH-1:0] out_868;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_868 (
            .a(out_867),
            .b(out_565),
            .outp(out_868)
        );        
        

        logic [WIDTH-1:0] out_869;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_869 (
            .a(out_866),
            .b(out_868),
            .outp(out_869)
        );        
        

        logic [WIDTH-1:0] out_870;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_870 (
            .in(out_869),
            .outp(out_870)
        );
        

        logic [WIDTH-1:0] out_871;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_871 (
            .a(out_865),
            .b(out_870),
            .outp(out_871)
        );        
        

        logic [WIDTH-1:0] out_872;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_872 (
            .a(out_863),
            .b(out_862),
            .outp(out_872)
        );        
        

        logic [WIDTH-1:0] out_873;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_873 (
            .a(out_869),
            .b(out_872),
            .outp(out_873)
        );        
        

        logic [WIDTH-1:0] out_874;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_874 (
            .in(out_861),
            .outp(out_874)
        );
        

        logic [WIDTH-1:0] out_875;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_875 (
            .a(out_873),
            .b(out_874),
            .outp(out_875)
        );        
        

        logic [WIDTH-1:0] out_876;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_876 (
            .a(out_871),
            .b(out_875),
            .outp(out_876)
        );        
        

        logic [WIDTH-1:0] out_877;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.813008)
        ) inst_877 (
            .outp(out_877)
        );
        

        logic [WIDTH-1:0] out_878;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_878 (
            .a(out_13),
            .b(out_877),
            .outp(out_878)
        );        
        

        logic [WIDTH-1:0] out_879;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.188)
        ) inst_879 (
            .outp(out_879)
        );
        

        logic [WIDTH-1:0] out_880;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_880 (
            .a(out_878),
            .b(out_879),
            .outp(out_880)
        );        
        

        logic [WIDTH-1:0] out_881;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_881 (
            .a(out_3),
            .b(out_880),
            .outp(out_881)
        );        
        

        logic [WIDTH-1:0] out_882;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0706995)
        ) inst_882 (
            .outp(out_882)
        );
        

        logic [WIDTH-1:0] out_883;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.60163)
        ) inst_883 (
            .outp(out_883)
        );
        

        logic [WIDTH-1:0] out_884;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_884 (
            .a(out_13),
            .b(out_883),
            .outp(out_884)
        );        
        

        logic [WIDTH-1:0] out_885;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_885 (
            .a(out_882),
            .b(out_884),
            .outp(out_885)
        );        
        

        logic [WIDTH-1:0] out_886;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_886 (
            .a(out_1),
            .b(out_123),
            .outp(out_886)
        );        
        

        logic [WIDTH-1:0] out_887;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_887 (
            .a(out_885),
            .b(out_886),
            .outp(out_887)
        );        
        

        logic [WIDTH-1:0] out_888;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_888 (
            .in(out_887),
            .outp(out_888)
        );
        

        logic [WIDTH-1:0] out_889;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_889 (
            .a(out_881),
            .b(out_888),
            .outp(out_889)
        );        
        

        logic [WIDTH-1:0] out_890;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.41463)
        ) inst_890 (
            .outp(out_890)
        );
        

        logic [WIDTH-1:0] out_891;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_891 (
            .a(out_13),
            .b(out_890),
            .outp(out_891)
        );        
        

        logic [WIDTH-1:0] out_892;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.9037)
        ) inst_892 (
            .outp(out_892)
        );
        

        logic [WIDTH-1:0] out_893;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_893 (
            .a(out_891),
            .b(out_892),
            .outp(out_893)
        );        
        

        logic [WIDTH-1:0] out_894;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_894 (
            .a(out_1),
            .b(out_552),
            .outp(out_894)
        );        
        

        logic [WIDTH-1:0] out_895;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_895 (
            .a(out_893),
            .b(out_894),
            .outp(out_895)
        );        
        

        logic [WIDTH-1:0] out_896;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_896 (
            .a(out_889),
            .b(out_895),
            .outp(out_896)
        );        
        

        logic [WIDTH-1:0] out_897;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_897 (
            .a(out_876),
            .b(out_896),
            .outp(out_897)
        );        
        

        logic [WIDTH-1:0] out_898;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.9037)
        ) inst_898 (
            .outp(out_898)
        );
        

        logic [WIDTH-1:0] out_899;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_899 (
            .a(out_891),
            .b(out_898),
            .outp(out_899)
        );        
        

        logic [WIDTH-1:0] out_900;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_900 (
            .a(out_894),
            .b(out_899),
            .outp(out_900)
        );        
        

        logic [WIDTH-1:0] out_901;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0706992)
        ) inst_901 (
            .outp(out_901)
        );
        

        logic [WIDTH-1:0] out_902;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_902 (
            .a(out_901),
            .b(out_884),
            .outp(out_902)
        );        
        

        logic [WIDTH-1:0] out_903;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_903 (
            .a(out_902),
            .b(out_886),
            .outp(out_903)
        );        
        

        logic [WIDTH-1:0] out_904;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_904 (
            .a(out_900),
            .b(out_903),
            .outp(out_904)
        );        
        

        logic [WIDTH-1:0] out_905;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_905 (
            .a(out_880),
            .b(out_3),
            .outp(out_905)
        );        
        

        logic [WIDTH-1:0] out_906;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_906 (
            .a(out_904),
            .b(out_905),
            .outp(out_906)
        );        
        

        logic [WIDTH-1:0] out_907;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_907 (
            .a(out_897),
            .b(out_906),
            .outp(out_907)
        );        
        

        logic [WIDTH-1:0] out_908;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.728)
        ) inst_908 (
            .outp(out_908)
        );
        

        logic [WIDTH-1:0] out_909;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.19512)
        ) inst_909 (
            .outp(out_909)
        );
        

        logic [WIDTH-1:0] out_910;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_910 (
            .a(out_13),
            .b(out_909),
            .outp(out_910)
        );        
        

        logic [WIDTH-1:0] out_911;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_911 (
            .a(out_908),
            .b(out_910),
            .outp(out_911)
        );        
        

        logic [WIDTH-1:0] out_912;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_912 (
            .in(out_911),
            .outp(out_912)
        );
        

        logic [WIDTH-1:0] out_913;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.8053)
        ) inst_913 (
            .outp(out_913)
        );
        

        logic [WIDTH-1:0] out_914;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_914 (
            .a(out_913),
            .b(out_886),
            .outp(out_914)
        );        
        

        logic [WIDTH-1:0] out_915;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_915 (
            .a(out_912),
            .b(out_914),
            .outp(out_915)
        );        
        

        logic [WIDTH-1:0] out_916;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_916 (
            .a(out_910),
            .b(out_886),
            .outp(out_916)
        );        
        

        logic [WIDTH-1:0] out_917;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.171801)
        ) inst_917 (
            .outp(out_917)
        );
        

        logic [WIDTH-1:0] out_918;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_918 (
            .a(out_916),
            .b(out_917),
            .outp(out_918)
        );        
        

        logic [WIDTH-1:0] out_919;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_919 (
            .a(out_915),
            .b(out_918),
            .outp(out_919)
        );        
        

        logic [WIDTH-1:0] out_920;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_920 (
            .a(out_907),
            .b(out_919),
            .outp(out_920)
        );        
        

        logic [WIDTH-1:0] out_921;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_921 (
            .a(out_917),
            .b(out_916),
            .outp(out_921)
        );        
        

        logic [WIDTH-1:0] out_922;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_922 (
            .a(out_911),
            .b(out_921),
            .outp(out_922)
        );        
        

        logic [WIDTH-1:0] out_923;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_923 (
            .a(out_886),
            .b(out_913),
            .outp(out_923)
        );        
        

        logic [WIDTH-1:0] out_924;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_924 (
            .a(out_922),
            .b(out_923),
            .outp(out_924)
        );        
        

        logic [WIDTH-1:0] out_925;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_925 (
            .a(out_920),
            .b(out_924),
            .outp(out_925)
        );        
        

        logic [WIDTH-1:0] out_926;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.12)
        ) inst_926 (
            .outp(out_926)
        );
        

        logic [WIDTH-1:0] out_927;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.25203)
        ) inst_927 (
            .outp(out_927)
        );
        

        logic [WIDTH-1:0] out_928;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_928 (
            .a(out_13),
            .b(out_927),
            .outp(out_928)
        );        
        

        logic [WIDTH-1:0] out_929;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_929 (
            .a(out_926),
            .b(out_928),
            .outp(out_929)
        );        
        

        logic [WIDTH-1:0] out_930;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.1769)
        ) inst_930 (
            .outp(out_930)
        );
        

        logic [WIDTH-1:0] out_931;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_931 (
            .a(out_928),
            .b(out_930),
            .outp(out_931)
        );        
        

        logic [WIDTH-1:0] out_932;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_932 (
            .a(out_127),
            .b(out_931),
            .outp(out_932)
        );        
        

        logic [WIDTH-1:0] out_933;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_933 (
            .a(out_929),
            .b(out_932),
            .outp(out_933)
        );        
        

        logic [WIDTH-1:0] out_934;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8369)
        ) inst_934 (
            .outp(out_934)
        );
        

        logic [WIDTH-1:0] out_935;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_935 (
            .a(out_934),
            .b(out_127),
            .outp(out_935)
        );        
        

        logic [WIDTH-1:0] out_936;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_936 (
            .a(out_933),
            .b(out_935),
            .outp(out_936)
        );        
        

        logic [WIDTH-1:0] out_937;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_937 (
            .a(out_925),
            .b(out_936),
            .outp(out_937)
        );        
        

        logic [WIDTH-1:0] out_938;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_938 (
            .a(out_127),
            .b(out_934),
            .outp(out_938)
        );        
        

        logic [WIDTH-1:0] out_939;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_939 (
            .a(out_931),
            .b(out_127),
            .outp(out_939)
        );        
        

        logic [WIDTH-1:0] out_940;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_940 (
            .a(out_938),
            .b(out_939),
            .outp(out_940)
        );        
        

        logic [WIDTH-1:0] out_941;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_941 (
            .in(out_929),
            .outp(out_941)
        );
        

        logic [WIDTH-1:0] out_942;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_942 (
            .a(out_940),
            .b(out_941),
            .outp(out_942)
        );        
        

        logic [WIDTH-1:0] out_943;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_943 (
            .a(out_937),
            .b(out_942),
            .outp(out_943)
        );        
        

        logic [WIDTH-1:0] out_944;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_944 (
            .in(out_943),
            .outp(out_944)
        );
        

        logic [WIDTH-1:0] out_945;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_945 (
            .a(out_944),
            .b(out_25),
            .outp(out_945)
        );        
        

        logic [WIDTH-1:0] out_946;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_946 (
            .a(out_945),
            .b(out_29),
            .outp(out_946)
        );        
        

        logic [WIDTH-1:0] out_947;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.558)
        ) inst_947 (
            .outp(out_947)
        );
        

        logic [WIDTH-1:0] out_948;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_948 (
            .a(out_3),
            .b(out_947),
            .outp(out_948)
        );        
        

        logic [WIDTH-1:0] out_949;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_949 (
            .a(out_946),
            .b(out_948),
            .outp(out_949)
        );        
        

        logic [WIDTH-1:0] out_950;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.058)
        ) inst_950 (
            .outp(out_950)
        );
        

        logic [WIDTH-1:0] out_951;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_951 (
            .a(out_950),
            .b(out_3),
            .outp(out_951)
        );        
        

        logic [WIDTH-1:0] out_952;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_952 (
            .a(out_949),
            .b(out_951),
            .outp(out_952)
        );        
        

        logic [WIDTH-1:0] out_953;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_953 (
            .a(out_859),
            .b(out_952),
            .outp(out_953)
        );        
        

        logic [WIDTH-1:0] out_954;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.683)
        ) inst_954 (
            .outp(out_954)
        );
        

        logic [WIDTH-1:0] out_955;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_955 (
            .a(out_3),
            .b(out_954),
            .outp(out_955)
        );        
        

        logic [WIDTH-1:0] out_956;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_956 (
            .in(out_955),
            .outp(out_956)
        );
        

        logic [WIDTH-1:0] out_957;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_957 (
            .a(out_16),
            .b(out_956),
            .outp(out_957)
        );        
        

        logic [WIDTH-1:0] out_958;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_958 (
            .in(out_957),
            .outp(out_958)
        );
        

        logic [WIDTH-1:0] out_959;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_959 (
            .a(out_9),
            .b(out_958),
            .outp(out_959)
        );        
        

        logic [WIDTH-1:0] out_960;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_960 (
            .a(out_958),
            .b(out_21),
            .outp(out_960)
        );        
        

        logic [WIDTH-1:0] out_961;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_961 (
            .a(out_959),
            .b(out_960),
            .outp(out_961)
        );        
        

        logic [WIDTH-1:0] out_962;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_962 (
            .a(out_953),
            .b(out_961),
            .outp(out_962)
        );        
        

        logic [WIDTH-1:0] out_963;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.033)
        ) inst_963 (
            .outp(out_963)
        );
        

        logic [WIDTH-1:0] out_964;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_964 (
            .a(out_3),
            .b(out_963),
            .outp(out_964)
        );        
        

        logic [WIDTH-1:0] out_965;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_965 (
            .in(out_964),
            .outp(out_965)
        );
        

        logic [WIDTH-1:0] out_966;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_966 (
            .a(out_16),
            .b(out_965),
            .outp(out_966)
        );        
        

        logic [WIDTH-1:0] out_967;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_967 (
            .in(out_966),
            .outp(out_967)
        );
        

        logic [WIDTH-1:0] out_968;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_968 (
            .a(out_9),
            .b(out_967),
            .outp(out_968)
        );        
        

        logic [WIDTH-1:0] out_969;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_969 (
            .a(out_967),
            .b(out_21),
            .outp(out_969)
        );        
        

        logic [WIDTH-1:0] out_970;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_970 (
            .a(out_968),
            .b(out_969),
            .outp(out_970)
        );        
        

        logic [WIDTH-1:0] out_971;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_971 (
            .a(out_962),
            .b(out_970),
            .outp(out_971)
        );        
        

        logic [WIDTH-1:0] out_972;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.233)
        ) inst_972 (
            .outp(out_972)
        );
        

        logic [WIDTH-1:0] out_973;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_973 (
            .a(out_3),
            .b(out_972),
            .outp(out_973)
        );        
        

        logic [WIDTH-1:0] out_974;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.133)
        ) inst_974 (
            .outp(out_974)
        );
        

        logic [WIDTH-1:0] out_975;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_975 (
            .a(out_974),
            .b(out_3),
            .outp(out_975)
        );        
        

        logic [WIDTH-1:0] out_976;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_976 (
            .a(out_973),
            .b(out_975),
            .outp(out_976)
        );        
        

        logic [WIDTH-1:0] out_977;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_977 (
            .a(out_976),
            .b(out_25),
            .outp(out_977)
        );        
        

        logic [WIDTH-1:0] out_978;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_978 (
            .a(out_977),
            .b(out_29),
            .outp(out_978)
        );        
        

        logic [WIDTH-1:0] out_979;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_979 (
            .a(out_971),
            .b(out_978),
            .outp(out_979)
        );        
        

        logic [WIDTH-1:0] out_980;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_980 (
            .a(out_52),
            .b(out_233),
            .outp(out_980)
        );        
        

        logic [WIDTH-1:0] out_981;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.408)
        ) inst_981 (
            .outp(out_981)
        );
        

        logic [WIDTH-1:0] out_982;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_982 (
            .a(out_3),
            .b(out_981),
            .outp(out_982)
        );        
        

        logic [WIDTH-1:0] out_983;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_983 (
            .a(out_980),
            .b(out_982),
            .outp(out_983)
        );        
        

        logic [WIDTH-1:0] out_984;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.233)
        ) inst_984 (
            .outp(out_984)
        );
        

        logic [WIDTH-1:0] out_985;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_985 (
            .a(out_984),
            .b(out_3),
            .outp(out_985)
        );        
        

        logic [WIDTH-1:0] out_986;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_986 (
            .a(out_983),
            .b(out_985),
            .outp(out_986)
        );        
        

        logic [WIDTH-1:0] out_987;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_987 (
            .a(out_979),
            .b(out_986),
            .outp(out_987)
        );        
        

        logic [WIDTH-1:0] out_988;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_988 (
            .a(out_982),
            .b(out_985),
            .outp(out_988)
        );        
        

        logic [WIDTH-1:0] out_989;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_989 (
            .a(out_988),
            .b(out_77),
            .outp(out_989)
        );        
        

        logic [WIDTH-1:0] out_990;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_990 (
            .a(out_989),
            .b(out_29),
            .outp(out_990)
        );        
        

        logic [WIDTH-1:0] out_991;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_991 (
            .a(out_987),
            .b(out_990),
            .outp(out_991)
        );        
        

        logic [WIDTH-1:0] out_992;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.133)
        ) inst_992 (
            .outp(out_992)
        );
        

        logic [WIDTH-1:0] out_993;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_993 (
            .a(out_3),
            .b(out_992),
            .outp(out_993)
        );        
        

        logic [WIDTH-1:0] out_994;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.408)
        ) inst_994 (
            .outp(out_994)
        );
        

        logic [WIDTH-1:0] out_995;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_995 (
            .a(out_994),
            .b(out_3),
            .outp(out_995)
        );        
        

        logic [WIDTH-1:0] out_996;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_996 (
            .a(out_993),
            .b(out_995),
            .outp(out_996)
        );        
        

        logic [WIDTH-1:0] out_997;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_997 (
            .in(out_982),
            .outp(out_997)
        );
        

        logic [WIDTH-1:0] out_998;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_998 (
            .a(out_16),
            .b(out_997),
            .outp(out_998)
        );        
        

        logic [WIDTH-1:0] out_999;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_999 (
            .in(out_998),
            .outp(out_999)
        );
        

        logic [WIDTH-1:0] out_1000;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1000 (
            .a(out_9),
            .b(out_999),
            .outp(out_1000)
        );        
        

        logic [WIDTH-1:0] out_1001;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1001 (
            .a(out_996),
            .b(out_1000),
            .outp(out_1001)
        );        
        

        logic [WIDTH-1:0] out_1002;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1002 (
            .a(out_999),
            .b(out_21),
            .outp(out_1002)
        );        
        

        logic [WIDTH-1:0] out_1003;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1003 (
            .a(out_1001),
            .b(out_1002),
            .outp(out_1003)
        );        
        

        logic [WIDTH-1:0] out_1004;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1004 (
            .a(out_1003),
            .b(out_25),
            .outp(out_1004)
        );        
        

        logic [WIDTH-1:0] out_1005;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1005 (
            .a(out_1004),
            .b(out_29),
            .outp(out_1005)
        );        
        

        logic [WIDTH-1:0] out_1006;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1006 (
            .a(out_991),
            .b(out_1005),
            .outp(out_1006)
        );        
        

        logic [WIDTH-1:0] out_1007;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.685)
        ) inst_1007 (
            .outp(out_1007)
        );
        

        logic [WIDTH-1:0] out_1008;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1008 (
            .a(out_1007),
            .b(out_152),
            .outp(out_1008)
        );        
        

        logic [WIDTH-1:0] out_1009;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1009 (
            .in(out_1008),
            .outp(out_1009)
        );
        

        logic [WIDTH-1:0] out_1010;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.82927)
        ) inst_1010 (
            .outp(out_1010)
        );
        

        logic [WIDTH-1:0] out_1011;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1011 (
            .a(out_13),
            .b(out_1010),
            .outp(out_1011)
        );        
        

        logic [WIDTH-1:0] out_1012;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5769)
        ) inst_1012 (
            .outp(out_1012)
        );
        

        logic [WIDTH-1:0] out_1013;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1013 (
            .a(out_1011),
            .b(out_1012),
            .outp(out_1013)
        );        
        

        logic [WIDTH-1:0] out_1014;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1014 (
            .a(out_127),
            .b(out_1013),
            .outp(out_1014)
        );        
        

        logic [WIDTH-1:0] out_1015;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1015 (
            .a(out_1009),
            .b(out_1014),
            .outp(out_1015)
        );        
        

        logic [WIDTH-1:0] out_1016;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.64228)
        ) inst_1016 (
            .outp(out_1016)
        );
        

        logic [WIDTH-1:0] out_1017;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1017 (
            .a(out_13),
            .b(out_1016),
            .outp(out_1017)
        );        
        

        logic [WIDTH-1:0] out_1018;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2069)
        ) inst_1018 (
            .outp(out_1018)
        );
        

        logic [WIDTH-1:0] out_1019;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1019 (
            .a(out_1017),
            .b(out_1018),
            .outp(out_1019)
        );        
        

        logic [WIDTH-1:0] out_1020;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1020 (
            .a(out_1019),
            .b(out_127),
            .outp(out_1020)
        );        
        

        logic [WIDTH-1:0] out_1021;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1021 (
            .a(out_1015),
            .b(out_1020),
            .outp(out_1021)
        );        
        

        logic [WIDTH-1:0] out_1022;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1022 (
            .a(out_1006),
            .b(out_1021),
            .outp(out_1022)
        );        
        

        logic [WIDTH-1:0] out_1023;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1023 (
            .a(out_127),
            .b(out_1019),
            .outp(out_1023)
        );        
        

        logic [WIDTH-1:0] out_1024;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1024 (
            .a(out_1008),
            .b(out_1023),
            .outp(out_1024)
        );        
        

        logic [WIDTH-1:0] out_1025;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1025 (
            .a(out_1013),
            .b(out_127),
            .outp(out_1025)
        );        
        

        logic [WIDTH-1:0] out_1026;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1026 (
            .a(out_1024),
            .b(out_1025),
            .outp(out_1026)
        );        
        

        logic [WIDTH-1:0] out_1027;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1027 (
            .a(out_1022),
            .b(out_1026),
            .outp(out_1027)
        );        
        

        logic [WIDTH-1:0] out_1028;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.083)
        ) inst_1028 (
            .outp(out_1028)
        );
        

        logic [WIDTH-1:0] out_1029;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1029 (
            .a(out_1028),
            .b(out_3),
            .outp(out_1029)
        );        
        

        logic [WIDTH-1:0] out_1030;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.65)
        ) inst_1030 (
            .outp(out_1030)
        );
        

        logic [WIDTH-1:0] out_1031;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1031 (
            .a(out_1030),
            .b(out_14),
            .outp(out_1031)
        );        
        

        logic [WIDTH-1:0] out_1032;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1032 (
            .a(out_1029),
            .b(out_1031),
            .outp(out_1032)
        );        
        

        logic [WIDTH-1:0] out_1033;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.95)
        ) inst_1033 (
            .outp(out_1033)
        );
        

        logic [WIDTH-1:0] out_1034;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1034 (
            .a(out_1033),
            .b(out_14),
            .outp(out_1034)
        );        
        

        logic [WIDTH-1:0] out_1035;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1035 (
            .in(out_1034),
            .outp(out_1035)
        );
        

        logic [WIDTH-1:0] out_1036;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1036 (
            .a(out_1032),
            .b(out_1035),
            .outp(out_1036)
        );        
        

        logic [WIDTH-1:0] out_1037;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.733)
        ) inst_1037 (
            .outp(out_1037)
        );
        

        logic [WIDTH-1:0] out_1038;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1038 (
            .a(out_3),
            .b(out_1037),
            .outp(out_1038)
        );        
        

        logic [WIDTH-1:0] out_1039;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1039 (
            .a(out_1036),
            .b(out_1038),
            .outp(out_1039)
        );        
        

        logic [WIDTH-1:0] out_1040;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.95)
        ) inst_1040 (
            .outp(out_1040)
        );
        

        logic [WIDTH-1:0] out_1041;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1041 (
            .a(out_1040),
            .b(out_14),
            .outp(out_1041)
        );        
        

        logic [WIDTH-1:0] out_1042;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1042 (
            .in(out_1041),
            .outp(out_1042)
        );
        

        logic [WIDTH-1:0] out_1043;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.508)
        ) inst_1043 (
            .outp(out_1043)
        );
        

        logic [WIDTH-1:0] out_1044;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1044 (
            .a(out_3),
            .b(out_1043),
            .outp(out_1044)
        );        
        

        logic [WIDTH-1:0] out_1045;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1045 (
            .in(out_1044),
            .outp(out_1045)
        );
        

        logic [WIDTH-1:0] out_1046;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1046 (
            .a(out_1042),
            .b(out_1045),
            .outp(out_1046)
        );        
        

        logic [WIDTH-1:0] out_1047;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1047 (
            .in(out_1046),
            .outp(out_1047)
        );
        

        logic [WIDTH-1:0] out_1048;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1048 (
            .a(out_460),
            .b(out_1047),
            .outp(out_1048)
        );        
        

        logic [WIDTH-1:0] out_1049;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1049 (
            .a(out_1047),
            .b(out_9),
            .outp(out_1049)
        );        
        

        logic [WIDTH-1:0] out_1050;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1050 (
            .a(out_1048),
            .b(out_1049),
            .outp(out_1050)
        );        
        

        logic [WIDTH-1:0] out_1051;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.258)
        ) inst_1051 (
            .outp(out_1051)
        );
        

        logic [WIDTH-1:0] out_1052;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1052 (
            .a(out_3),
            .b(out_1051),
            .outp(out_1052)
        );        
        

        logic [WIDTH-1:0] out_1053;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1053 (
            .in(out_1052),
            .outp(out_1053)
        );
        

        logic [WIDTH-1:0] out_1054;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1054 (
            .a(out_1042),
            .b(out_1053),
            .outp(out_1054)
        );        
        

        logic [WIDTH-1:0] out_1055;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1055 (
            .in(out_1054),
            .outp(out_1055)
        );
        

        logic [WIDTH-1:0] out_1056;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1056 (
            .a(out_460),
            .b(out_1055),
            .outp(out_1056)
        );        
        

        logic [WIDTH-1:0] out_1057;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1057 (
            .a(out_1055),
            .b(out_9),
            .outp(out_1057)
        );        
        

        logic [WIDTH-1:0] out_1058;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1058 (
            .a(out_1056),
            .b(out_1057),
            .outp(out_1058)
        );        
        

        logic [WIDTH-1:0] out_1059;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1059 (
            .a(out_1050),
            .b(out_1058),
            .outp(out_1059)
        );        
        

        logic [WIDTH-1:0] out_1060;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1060 (
            .a(out_1039),
            .b(out_1059),
            .outp(out_1060)
        );        
        

        logic [WIDTH-1:0] out_1061;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1061 (
            .a(out_1027),
            .b(out_1060),
            .outp(out_1061)
        );        
        

        logic [WIDTH-1:0] out_1062;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.975)
        ) inst_1062 (
            .outp(out_1062)
        );
        

        logic [WIDTH-1:0] out_1063;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1063 (
            .a(out_1062),
            .b(out_14),
            .outp(out_1063)
        );        
        

        logic [WIDTH-1:0] out_1064;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1064 (
            .a(out_29),
            .b(out_1063),
            .outp(out_1064)
        );        
        

        logic [WIDTH-1:0] out_1065;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.282999)
        ) inst_1065 (
            .outp(out_1065)
        );
        

        logic [WIDTH-1:0] out_1066;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1066 (
            .a(out_3),
            .b(out_1065),
            .outp(out_1066)
        );        
        

        logic [WIDTH-1:0] out_1067;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1067 (
            .a(out_1064),
            .b(out_1066),
            .outp(out_1067)
        );        
        

        logic [WIDTH-1:0] out_1068;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.182999)
        ) inst_1068 (
            .outp(out_1068)
        );
        

        logic [WIDTH-1:0] out_1069;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1069 (
            .a(out_1068),
            .b(out_3),
            .outp(out_1069)
        );        
        

        logic [WIDTH-1:0] out_1070;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1070 (
            .a(out_1067),
            .b(out_1069),
            .outp(out_1070)
        );        
        

        logic [WIDTH-1:0] out_1071;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1071 (
            .a(out_1061),
            .b(out_1070),
            .outp(out_1071)
        );        
        

        logic [WIDTH-1:0] out_1072;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1072 (
            .a(out_52),
            .b(out_29),
            .outp(out_1072)
        );        
        

        logic [WIDTH-1:0] out_1073;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.167001)
        ) inst_1073 (
            .outp(out_1073)
        );
        

        logic [WIDTH-1:0] out_1074;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1074 (
            .a(out_1073),
            .b(out_3),
            .outp(out_1074)
        );        
        

        logic [WIDTH-1:0] out_1075;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1075 (
            .a(out_1072),
            .b(out_1074),
            .outp(out_1075)
        );        
        

        logic [WIDTH-1:0] out_1076;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.267001)
        ) inst_1076 (
            .outp(out_1076)
        );
        

        logic [WIDTH-1:0] out_1077;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1077 (
            .a(out_1076),
            .b(out_3),
            .outp(out_1077)
        );        
        

        logic [WIDTH-1:0] out_1078;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1078 (
            .in(out_1077),
            .outp(out_1078)
        );
        

        logic [WIDTH-1:0] out_1079;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1079 (
            .a(out_1075),
            .b(out_1078),
            .outp(out_1079)
        );        
        

        logic [WIDTH-1:0] out_1080;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1080 (
            .a(out_1071),
            .b(out_1079),
            .outp(out_1080)
        );        
        

        logic [WIDTH-1:0] out_1081;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1081 (
            .a(out_52),
            .b(out_1066),
            .outp(out_1081)
        );        
        

        logic [WIDTH-1:0] out_1082;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1082 (
            .a(out_1081),
            .b(out_1078),
            .outp(out_1082)
        );        
        

        logic [WIDTH-1:0] out_1083;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1083 (
            .in(out_1063),
            .outp(out_1083)
        );
        

        logic [WIDTH-1:0] out_1084;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1084 (
            .a(out_1082),
            .b(out_1083),
            .outp(out_1084)
        );        
        

        logic [WIDTH-1:0] out_1085;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.00799847)
        ) inst_1085 (
            .outp(out_1085)
        );
        

        logic [WIDTH-1:0] out_1086;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1086 (
            .a(out_3),
            .b(out_1085),
            .outp(out_1086)
        );        
        

        logic [WIDTH-1:0] out_1087;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1087 (
            .in(out_1086),
            .outp(out_1087)
        );
        

        logic [WIDTH-1:0] out_1088;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1088 (
            .a(out_16),
            .b(out_1087),
            .outp(out_1088)
        );        
        

        logic [WIDTH-1:0] out_1089;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1089 (
            .in(out_1088),
            .outp(out_1089)
        );
        

        logic [WIDTH-1:0] out_1090;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1090 (
            .a(out_9),
            .b(out_1089),
            .outp(out_1090)
        );        
        

        logic [WIDTH-1:0] out_1091;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1091 (
            .a(out_1084),
            .b(out_1090),
            .outp(out_1091)
        );        
        

        logic [WIDTH-1:0] out_1092;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1092 (
            .a(out_1089),
            .b(out_21),
            .outp(out_1092)
        );        
        

        logic [WIDTH-1:0] out_1093;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1093 (
            .a(out_1091),
            .b(out_1092),
            .outp(out_1093)
        );        
        

        logic [WIDTH-1:0] out_1094;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1094 (
            .a(out_1080),
            .b(out_1093),
            .outp(out_1094)
        );        
        

        logic [WIDTH-1:0] out_1095;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.23565)
        ) inst_1095 (
            .outp(out_1095)
        );
        

        logic [WIDTH-1:0] out_1096;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1096 (
            .a(out_1095),
            .b(out_131),
            .outp(out_1096)
        );        
        

        logic [WIDTH-1:0] out_1097;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1097 (
            .a(out_127),
            .b(out_1096),
            .outp(out_1097)
        );        
        

        logic [WIDTH-1:0] out_1098;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.81065)
        ) inst_1098 (
            .outp(out_1098)
        );
        

        logic [WIDTH-1:0] out_1099;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1099 (
            .a(out_1098),
            .b(out_124),
            .outp(out_1099)
        );        
        

        logic [WIDTH-1:0] out_1100;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1100 (
            .a(out_1099),
            .b(out_127),
            .outp(out_1100)
        );        
        

        logic [WIDTH-1:0] out_1101;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1101 (
            .a(out_1097),
            .b(out_1100),
            .outp(out_1101)
        );        
        

        logic [WIDTH-1:0] out_1102;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1102 (
            .a(out_1101),
            .b(out_154),
            .outp(out_1102)
        );        
        

        logic [WIDTH-1:0] out_1103;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1103 (
            .a(out_1094),
            .b(out_1102),
            .outp(out_1103)
        );        
        

        logic [WIDTH-1:0] out_1104;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1104 (
            .a(out_127),
            .b(out_1099),
            .outp(out_1104)
        );        
        

        logic [WIDTH-1:0] out_1105;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1105 (
            .a(out_1096),
            .b(out_127),
            .outp(out_1105)
        );        
        

        logic [WIDTH-1:0] out_1106;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1106 (
            .a(out_1104),
            .b(out_1105),
            .outp(out_1106)
        );        
        

        logic [WIDTH-1:0] out_1107;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1107 (
            .a(out_1106),
            .b(out_153),
            .outp(out_1107)
        );        
        

        logic [WIDTH-1:0] out_1108;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1108 (
            .a(out_1103),
            .b(out_1107),
            .outp(out_1108)
        );        
        

        logic [WIDTH-1:0] out_1109;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.18065)
        ) inst_1109 (
            .outp(out_1109)
        );
        

        logic [WIDTH-1:0] out_1110;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1110 (
            .a(out_1109),
            .b(out_131),
            .outp(out_1110)
        );        
        

        logic [WIDTH-1:0] out_1111;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1111 (
            .a(out_1110),
            .b(out_127),
            .outp(out_1111)
        );        
        

        logic [WIDTH-1:0] out_1112;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1112 (
            .a(out_1104),
            .b(out_1111),
            .outp(out_1112)
        );        
        

        logic [WIDTH-1:0] out_1113;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1113 (
            .a(out_1112),
            .b(out_138),
            .outp(out_1113)
        );        
        

        logic [WIDTH-1:0] out_1114;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1114 (
            .a(out_1108),
            .b(out_1113),
            .outp(out_1114)
        );        
        

        logic [WIDTH-1:0] out_1115;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1115 (
            .a(out_127),
            .b(out_1110),
            .outp(out_1115)
        );        
        

        logic [WIDTH-1:0] out_1116;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1116 (
            .a(out_1100),
            .b(out_1115),
            .outp(out_1116)
        );        
        

        logic [WIDTH-1:0] out_1117;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1117 (
            .a(out_1116),
            .b(out_139),
            .outp(out_1117)
        );        
        

        logic [WIDTH-1:0] out_1118;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1118 (
            .a(out_1114),
            .b(out_1117),
            .outp(out_1118)
        );        
        

        logic [WIDTH-1:0] out_1119;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.96935)
        ) inst_1119 (
            .outp(out_1119)
        );
        

        logic [WIDTH-1:0] out_1120;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1120 (
            .a(out_1119),
            .b(out_131),
            .outp(out_1120)
        );        
        

        logic [WIDTH-1:0] out_1121;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1121 (
            .a(out_1120),
            .b(out_127),
            .outp(out_1121)
        );        
        

        logic [WIDTH-1:0] out_1122;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1122 (
            .in(out_1121),
            .outp(out_1122)
        );
        

        logic [WIDTH-1:0] out_1123;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.54435)
        ) inst_1123 (
            .outp(out_1123)
        );
        

        logic [WIDTH-1:0] out_1124;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1124 (
            .a(out_1123),
            .b(out_124),
            .outp(out_1124)
        );        
        

        logic [WIDTH-1:0] out_1125;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1125 (
            .a(out_1124),
            .b(out_127),
            .outp(out_1125)
        );        
        

        logic [WIDTH-1:0] out_1126;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1126 (
            .a(out_1122),
            .b(out_1125),
            .outp(out_1126)
        );        
        

        logic [WIDTH-1:0] out_1127;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1127 (
            .a(out_1126),
            .b(out_154),
            .outp(out_1127)
        );        
        

        logic [WIDTH-1:0] out_1128;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1128 (
            .a(out_1118),
            .b(out_1127),
            .outp(out_1128)
        );        
        

        logic [WIDTH-1:0] out_1129;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1129 (
            .in(out_1125),
            .outp(out_1129)
        );
        

        logic [WIDTH-1:0] out_1130;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1130 (
            .a(out_1121),
            .b(out_1129),
            .outp(out_1130)
        );        
        

        logic [WIDTH-1:0] out_1131;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1131 (
            .a(out_1130),
            .b(out_153),
            .outp(out_1131)
        );        
        

        logic [WIDTH-1:0] out_1132;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1132 (
            .a(out_1128),
            .b(out_1131),
            .outp(out_1132)
        );        
        

        logic [WIDTH-1:0] out_1133;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.91435)
        ) inst_1133 (
            .outp(out_1133)
        );
        

        logic [WIDTH-1:0] out_1134;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1134 (
            .a(out_1133),
            .b(out_131),
            .outp(out_1134)
        );        
        

        logic [WIDTH-1:0] out_1135;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1135 (
            .a(out_1134),
            .b(out_127),
            .outp(out_1135)
        );        
        

        logic [WIDTH-1:0] out_1136;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1136 (
            .a(out_1129),
            .b(out_1135),
            .outp(out_1136)
        );        
        

        logic [WIDTH-1:0] out_1137;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1137 (
            .a(out_1136),
            .b(out_138),
            .outp(out_1137)
        );        
        

        logic [WIDTH-1:0] out_1138;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1138 (
            .a(out_1132),
            .b(out_1137),
            .outp(out_1138)
        );        
        

        logic [WIDTH-1:0] out_1139;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1139 (
            .in(out_1135),
            .outp(out_1139)
        );
        

        logic [WIDTH-1:0] out_1140;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1140 (
            .a(out_1125),
            .b(out_1139),
            .outp(out_1140)
        );        
        

        logic [WIDTH-1:0] out_1141;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1141 (
            .a(out_1140),
            .b(out_139),
            .outp(out_1141)
        );        
        

        logic [WIDTH-1:0] out_1142;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1142 (
            .a(out_1138),
            .b(out_1141),
            .outp(out_1142)
        );        
        

        logic [WIDTH-1:0] out_1143;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.96065)
        ) inst_1143 (
            .outp(out_1143)
        );
        

        logic [WIDTH-1:0] out_1144;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1144 (
            .a(out_1143),
            .b(out_131),
            .outp(out_1144)
        );        
        

        logic [WIDTH-1:0] out_1145;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1145 (
            .a(out_127),
            .b(out_1144),
            .outp(out_1145)
        );        
        

        logic [WIDTH-1:0] out_1146;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1146 (
            .a(out_1145),
            .b(out_128),
            .outp(out_1146)
        );        
        

        logic [WIDTH-1:0] out_1147;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1147 (
            .a(out_1146),
            .b(out_154),
            .outp(out_1147)
        );        
        

        logic [WIDTH-1:0] out_1148;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1148 (
            .a(out_1142),
            .b(out_1147),
            .outp(out_1148)
        );        
        

        logic [WIDTH-1:0] out_1149;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.53565)
        ) inst_1149 (
            .outp(out_1149)
        );
        

        logic [WIDTH-1:0] out_1150;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1150 (
            .a(out_1149),
            .b(out_124),
            .outp(out_1150)
        );        
        

        logic [WIDTH-1:0] out_1151;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1151 (
            .a(out_127),
            .b(out_1150),
            .outp(out_1151)
        );        
        

        logic [WIDTH-1:0] out_1152;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1152 (
            .a(out_1144),
            .b(out_127),
            .outp(out_1152)
        );        
        

        logic [WIDTH-1:0] out_1153;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1153 (
            .a(out_1151),
            .b(out_1152),
            .outp(out_1153)
        );        
        

        logic [WIDTH-1:0] out_1154;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1154 (
            .a(out_1153),
            .b(out_153),
            .outp(out_1154)
        );        
        

        logic [WIDTH-1:0] out_1155;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1155 (
            .a(out_1148),
            .b(out_1154),
            .outp(out_1155)
        );        
        

        logic [WIDTH-1:0] out_1156;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1156 (
            .a(out_132),
            .b(out_127),
            .outp(out_1156)
        );        
        

        logic [WIDTH-1:0] out_1157;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1157 (
            .a(out_1151),
            .b(out_1156),
            .outp(out_1157)
        );        
        

        logic [WIDTH-1:0] out_1158;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1158 (
            .a(out_1157),
            .b(out_138),
            .outp(out_1158)
        );        
        

        logic [WIDTH-1:0] out_1159;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1159 (
            .a(out_1155),
            .b(out_1158),
            .outp(out_1159)
        );        
        

        logic [WIDTH-1:0] out_1160;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.63)
        ) inst_1160 (
            .outp(out_1160)
        );
        

        logic [WIDTH-1:0] out_1161;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1161 (
            .a(out_1160),
            .b(out_137),
            .outp(out_1161)
        );        
        

        logic [WIDTH-1:0] out_1162;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1162 (
            .a(out_1023),
            .b(out_1161),
            .outp(out_1162)
        );        
        

        logic [WIDTH-1:0] out_1163;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5219)
        ) inst_1163 (
            .outp(out_1163)
        );
        

        logic [WIDTH-1:0] out_1164;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1164 (
            .a(out_1011),
            .b(out_1163),
            .outp(out_1164)
        );        
        

        logic [WIDTH-1:0] out_1165;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1165 (
            .a(out_1164),
            .b(out_127),
            .outp(out_1165)
        );        
        

        logic [WIDTH-1:0] out_1166;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1166 (
            .a(out_1162),
            .b(out_1165),
            .outp(out_1166)
        );        
        

        logic [WIDTH-1:0] out_1167;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1167 (
            .a(out_1159),
            .b(out_1166),
            .outp(out_1167)
        );        
        

        logic [WIDTH-1:0] out_1168;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1168 (
            .a(out_127),
            .b(out_1164),
            .outp(out_1168)
        );        
        

        logic [WIDTH-1:0] out_1169;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1169 (
            .a(out_1020),
            .b(out_1168),
            .outp(out_1169)
        );        
        

        logic [WIDTH-1:0] out_1170;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1170 (
            .in(out_1161),
            .outp(out_1170)
        );
        

        logic [WIDTH-1:0] out_1171;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1171 (
            .a(out_1169),
            .b(out_1170),
            .outp(out_1171)
        );        
        

        logic [WIDTH-1:0] out_1172;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1172 (
            .a(out_1167),
            .b(out_1171),
            .outp(out_1172)
        );        
        

        logic [WIDTH-1:0] out_1173;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1173 (
            .a(out_1014),
            .b(out_154),
            .outp(out_1173)
        );        
        

        logic [WIDTH-1:0] out_1174;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1519)
        ) inst_1174 (
            .outp(out_1174)
        );
        

        logic [WIDTH-1:0] out_1175;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1175 (
            .a(out_1017),
            .b(out_1174),
            .outp(out_1175)
        );        
        

        logic [WIDTH-1:0] out_1176;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1176 (
            .a(out_1175),
            .b(out_127),
            .outp(out_1176)
        );        
        

        logic [WIDTH-1:0] out_1177;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1177 (
            .a(out_1173),
            .b(out_1176),
            .outp(out_1177)
        );        
        

        logic [WIDTH-1:0] out_1178;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1178 (
            .a(out_1172),
            .b(out_1177),
            .outp(out_1178)
        );        
        

        logic [WIDTH-1:0] out_1179;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1179 (
            .a(out_1025),
            .b(out_153),
            .outp(out_1179)
        );        
        

        logic [WIDTH-1:0] out_1180;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1180 (
            .a(out_127),
            .b(out_1175),
            .outp(out_1180)
        );        
        

        logic [WIDTH-1:0] out_1181;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1181 (
            .a(out_1179),
            .b(out_1180),
            .outp(out_1181)
        );        
        

        logic [WIDTH-1:0] out_1182;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1182 (
            .a(out_1178),
            .b(out_1181),
            .outp(out_1182)
        );        
        

        logic [WIDTH-1:0] out_1183;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1183 (
            .a(out_1165),
            .b(out_1180),
            .outp(out_1183)
        );        
        

        logic [WIDTH-1:0] out_1184;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1184 (
            .a(out_1183),
            .b(out_138),
            .outp(out_1184)
        );        
        

        logic [WIDTH-1:0] out_1185;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1185 (
            .a(out_1182),
            .b(out_1184),
            .outp(out_1185)
        );        
        

        logic [WIDTH-1:0] out_1186;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1186 (
            .a(out_1168),
            .b(out_1176),
            .outp(out_1186)
        );        
        

        logic [WIDTH-1:0] out_1187;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1187 (
            .a(out_1186),
            .b(out_139),
            .outp(out_1187)
        );        
        

        logic [WIDTH-1:0] out_1188;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1188 (
            .a(out_1185),
            .b(out_1187),
            .outp(out_1188)
        );        
        

        logic [WIDTH-1:0] out_1189;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.3131)
        ) inst_1189 (
            .outp(out_1189)
        );
        

        logic [WIDTH-1:0] out_1190;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1190 (
            .a(out_1189),
            .b(out_1011),
            .outp(out_1190)
        );        
        

        logic [WIDTH-1:0] out_1191;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1191 (
            .a(out_1190),
            .b(out_127),
            .outp(out_1191)
        );        
        

        logic [WIDTH-1:0] out_1192;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1192 (
            .in(out_1191),
            .outp(out_1192)
        );
        

        logic [WIDTH-1:0] out_1193;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1193 (
            .a(out_154),
            .b(out_1192),
            .outp(out_1193)
        );        
        

        logic [WIDTH-1:0] out_1194;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.8881)
        ) inst_1194 (
            .outp(out_1194)
        );
        

        logic [WIDTH-1:0] out_1195;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1195 (
            .a(out_1194),
            .b(out_1017),
            .outp(out_1195)
        );        
        

        logic [WIDTH-1:0] out_1196;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1196 (
            .a(out_1195),
            .b(out_127),
            .outp(out_1196)
        );        
        

        logic [WIDTH-1:0] out_1197;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1197 (
            .a(out_1193),
            .b(out_1196),
            .outp(out_1197)
        );        
        

        logic [WIDTH-1:0] out_1198;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1198 (
            .a(out_1188),
            .b(out_1197),
            .outp(out_1198)
        );        
        

        logic [WIDTH-1:0] out_1199;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1199 (
            .a(out_153),
            .b(out_1191),
            .outp(out_1199)
        );        
        

        logic [WIDTH-1:0] out_1200;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1200 (
            .in(out_1196),
            .outp(out_1200)
        );
        

        logic [WIDTH-1:0] out_1201;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1201 (
            .a(out_1199),
            .b(out_1200),
            .outp(out_1201)
        );        
        

        logic [WIDTH-1:0] out_1202;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1202 (
            .a(out_1198),
            .b(out_1201),
            .outp(out_1202)
        );        
        

        logic [WIDTH-1:0] out_1203;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1203 (
            .a(out_138),
            .b(out_1200),
            .outp(out_1203)
        );        
        

        logic [WIDTH-1:0] out_1204;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.2581)
        ) inst_1204 (
            .outp(out_1204)
        );
        

        logic [WIDTH-1:0] out_1205;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1205 (
            .a(out_1204),
            .b(out_1011),
            .outp(out_1205)
        );        
        

        logic [WIDTH-1:0] out_1206;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1206 (
            .a(out_1205),
            .b(out_127),
            .outp(out_1206)
        );        
        

        logic [WIDTH-1:0] out_1207;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1207 (
            .a(out_1203),
            .b(out_1206),
            .outp(out_1207)
        );        
        

        logic [WIDTH-1:0] out_1208;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1208 (
            .a(out_1202),
            .b(out_1207),
            .outp(out_1208)
        );        
        

        logic [WIDTH-1:0] out_1209;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1209 (
            .a(out_139),
            .b(out_1196),
            .outp(out_1209)
        );        
        

        logic [WIDTH-1:0] out_1210;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1210 (
            .in(out_1206),
            .outp(out_1210)
        );
        

        logic [WIDTH-1:0] out_1211;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1211 (
            .a(out_1209),
            .b(out_1210),
            .outp(out_1211)
        );        
        

        logic [WIDTH-1:0] out_1212;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1212 (
            .a(out_1208),
            .b(out_1211),
            .outp(out_1212)
        );        
        

        logic [WIDTH-1:0] out_1213;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1213 (
            .a(out_29),
            .b(out_1041),
            .outp(out_1213)
        );        
        

        logic [WIDTH-1:0] out_1214;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.683)
        ) inst_1214 (
            .outp(out_1214)
        );
        

        logic [WIDTH-1:0] out_1215;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1215 (
            .a(out_3),
            .b(out_1214),
            .outp(out_1215)
        );        
        

        logic [WIDTH-1:0] out_1216;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1216 (
            .a(out_1213),
            .b(out_1215),
            .outp(out_1216)
        );        
        

        logic [WIDTH-1:0] out_1217;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.583)
        ) inst_1217 (
            .outp(out_1217)
        );
        

        logic [WIDTH-1:0] out_1218;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1218 (
            .a(out_1217),
            .b(out_3),
            .outp(out_1218)
        );        
        

        logic [WIDTH-1:0] out_1219;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1219 (
            .a(out_1216),
            .b(out_1218),
            .outp(out_1219)
        );        
        

        logic [WIDTH-1:0] out_1220;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1220 (
            .a(out_1212),
            .b(out_1219),
            .outp(out_1220)
        );        
        

        logic [WIDTH-1:0] out_1221;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.433)
        ) inst_1221 (
            .outp(out_1221)
        );
        

        logic [WIDTH-1:0] out_1222;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1222 (
            .a(out_3),
            .b(out_1221),
            .outp(out_1222)
        );        
        

        logic [WIDTH-1:0] out_1223;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1223 (
            .a(out_1213),
            .b(out_1222),
            .outp(out_1223)
        );        
        

        logic [WIDTH-1:0] out_1224;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.333)
        ) inst_1224 (
            .outp(out_1224)
        );
        

        logic [WIDTH-1:0] out_1225;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1225 (
            .a(out_1224),
            .b(out_3),
            .outp(out_1225)
        );        
        

        logic [WIDTH-1:0] out_1226;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1226 (
            .a(out_1223),
            .b(out_1225),
            .outp(out_1226)
        );        
        

        logic [WIDTH-1:0] out_1227;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1227 (
            .a(out_1220),
            .b(out_1226),
            .outp(out_1227)
        );        
        

        logic [WIDTH-1:0] out_1228;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.775)
        ) inst_1228 (
            .outp(out_1228)
        );
        

        logic [WIDTH-1:0] out_1229;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1229 (
            .a(out_1228),
            .b(out_14),
            .outp(out_1229)
        );        
        

        logic [WIDTH-1:0] out_1230;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1230 (
            .a(out_29),
            .b(out_1229),
            .outp(out_1230)
        );        
        

        logic [WIDTH-1:0] out_1231;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1231 (
            .a(out_1230),
            .b(out_546),
            .outp(out_1231)
        );        
        

        logic [WIDTH-1:0] out_1232;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1232 (
            .a(out_1231),
            .b(out_1029),
            .outp(out_1232)
        );        
        

        logic [WIDTH-1:0] out_1233;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1233 (
            .a(out_1227),
            .b(out_1232),
            .outp(out_1233)
        );        
        

        logic [WIDTH-1:0] out_1234;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.65)
        ) inst_1234 (
            .outp(out_1234)
        );
        

        logic [WIDTH-1:0] out_1235;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1235 (
            .a(out_1234),
            .b(out_14),
            .outp(out_1235)
        );        
        

        logic [WIDTH-1:0] out_1236;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.498)
        ) inst_1236 (
            .outp(out_1236)
        );
        

        logic [WIDTH-1:0] out_1237;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1237 (
            .a(out_3),
            .b(out_1236),
            .outp(out_1237)
        );        
        

        logic [WIDTH-1:0] out_1238;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1238 (
            .a(out_1235),
            .b(out_1237),
            .outp(out_1238)
        );        
        

        logic [WIDTH-1:0] out_1239;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.398)
        ) inst_1239 (
            .outp(out_1239)
        );
        

        logic [WIDTH-1:0] out_1240;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1240 (
            .a(out_1239),
            .b(out_3),
            .outp(out_1240)
        );        
        

        logic [WIDTH-1:0] out_1241;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1241 (
            .a(out_1238),
            .b(out_1240),
            .outp(out_1241)
        );        
        

        logic [WIDTH-1:0] out_1242;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0)
        ) inst_1242 (
            .outp(out_1242)
        );
        

        logic [WIDTH-1:0] out_1243;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1243 (
            .a(out_1242),
            .b(out_14),
            .outp(out_1243)
        );        
        

        logic [WIDTH-1:0] out_1244;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1244 (
            .in(out_1243),
            .outp(out_1244)
        );
        

        logic [WIDTH-1:0] out_1245;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1245 (
            .a(out_1241),
            .b(out_1244),
            .outp(out_1245)
        );        
        

        logic [WIDTH-1:0] out_1246;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1246 (
            .a(out_1233),
            .b(out_1245),
            .outp(out_1246)
        );        
        

        logic [WIDTH-1:0] out_1247;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.248)
        ) inst_1247 (
            .outp(out_1247)
        );
        

        logic [WIDTH-1:0] out_1248;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1248 (
            .a(out_3),
            .b(out_1247),
            .outp(out_1248)
        );        
        

        logic [WIDTH-1:0] out_1249;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1249 (
            .a(out_1235),
            .b(out_1248),
            .outp(out_1249)
        );        
        

        logic [WIDTH-1:0] out_1250;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.148)
        ) inst_1250 (
            .outp(out_1250)
        );
        

        logic [WIDTH-1:0] out_1251;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1251 (
            .a(out_1250),
            .b(out_3),
            .outp(out_1251)
        );        
        

        logic [WIDTH-1:0] out_1252;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1252 (
            .a(out_1249),
            .b(out_1251),
            .outp(out_1252)
        );        
        

        logic [WIDTH-1:0] out_1253;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1253 (
            .a(out_1252),
            .b(out_1244),
            .outp(out_1253)
        );        
        

        logic [WIDTH-1:0] out_1254;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1254 (
            .a(out_1246),
            .b(out_1253),
            .outp(out_1254)
        );        
        

        logic [WIDTH-1:0] out_1255;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.475)
        ) inst_1255 (
            .outp(out_1255)
        );
        

        logic [WIDTH-1:0] out_1256;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1256 (
            .a(out_1255),
            .b(out_14),
            .outp(out_1256)
        );        
        

        logic [WIDTH-1:0] out_1257;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.998001)
        ) inst_1257 (
            .outp(out_1257)
        );
        

        logic [WIDTH-1:0] out_1258;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1258 (
            .a(out_3),
            .b(out_1257),
            .outp(out_1258)
        );        
        

        logic [WIDTH-1:0] out_1259;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1259 (
            .a(out_1256),
            .b(out_1258),
            .outp(out_1259)
        );        
        

        logic [WIDTH-1:0] out_1260;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.898001)
        ) inst_1260 (
            .outp(out_1260)
        );
        

        logic [WIDTH-1:0] out_1261;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1261 (
            .a(out_1260),
            .b(out_3),
            .outp(out_1261)
        );        
        

        logic [WIDTH-1:0] out_1262;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1262 (
            .a(out_1259),
            .b(out_1261),
            .outp(out_1262)
        );        
        

        logic [WIDTH-1:0] out_1263;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1263 (
            .a(out_1262),
            .b(out_1244),
            .outp(out_1263)
        );        
        

        logic [WIDTH-1:0] out_1264;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1264 (
            .a(out_1254),
            .b(out_1263),
            .outp(out_1264)
        );        
        

        logic [WIDTH-1:0] out_1265;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.65)
        ) inst_1265 (
            .outp(out_1265)
        );
        

        logic [WIDTH-1:0] out_1266;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1266 (
            .a(out_1265),
            .b(out_14),
            .outp(out_1266)
        );        
        

        logic [WIDTH-1:0] out_1267;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1267 (
            .in(out_1266),
            .outp(out_1267)
        );
        

        logic [WIDTH-1:0] out_1268;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1268 (
            .a(out_1261),
            .b(out_1267),
            .outp(out_1268)
        );        
        

        logic [WIDTH-1:0] out_1269;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.548)
        ) inst_1269 (
            .outp(out_1269)
        );
        

        logic [WIDTH-1:0] out_1270;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1270 (
            .a(out_3),
            .b(out_1269),
            .outp(out_1270)
        );        
        

        logic [WIDTH-1:0] out_1271;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1271 (
            .a(out_1268),
            .b(out_1270),
            .outp(out_1271)
        );        
        

        logic [WIDTH-1:0] out_1272;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1272 (
            .in(out_1235),
            .outp(out_1272)
        );
        

        logic [WIDTH-1:0] out_1273;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.323)
        ) inst_1273 (
            .outp(out_1273)
        );
        

        logic [WIDTH-1:0] out_1274;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1274 (
            .a(out_3),
            .b(out_1273),
            .outp(out_1274)
        );        
        

        logic [WIDTH-1:0] out_1275;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1275 (
            .in(out_1274),
            .outp(out_1275)
        );
        

        logic [WIDTH-1:0] out_1276;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1276 (
            .a(out_1272),
            .b(out_1275),
            .outp(out_1276)
        );        
        

        logic [WIDTH-1:0] out_1277;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1277 (
            .in(out_1276),
            .outp(out_1277)
        );
        

        logic [WIDTH-1:0] out_1278;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1278 (
            .a(out_460),
            .b(out_1277),
            .outp(out_1278)
        );        
        

        logic [WIDTH-1:0] out_1279;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1279 (
            .a(out_1277),
            .b(out_9),
            .outp(out_1279)
        );        
        

        logic [WIDTH-1:0] out_1280;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1280 (
            .a(out_1278),
            .b(out_1279),
            .outp(out_1280)
        );        
        

        logic [WIDTH-1:0] out_1281;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.073)
        ) inst_1281 (
            .outp(out_1281)
        );
        

        logic [WIDTH-1:0] out_1282;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1282 (
            .a(out_3),
            .b(out_1281),
            .outp(out_1282)
        );        
        

        logic [WIDTH-1:0] out_1283;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1283 (
            .in(out_1282),
            .outp(out_1283)
        );
        

        logic [WIDTH-1:0] out_1284;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1284 (
            .a(out_1272),
            .b(out_1283),
            .outp(out_1284)
        );        
        

        logic [WIDTH-1:0] out_1285;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1285 (
            .in(out_1284),
            .outp(out_1285)
        );
        

        logic [WIDTH-1:0] out_1286;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1286 (
            .a(out_460),
            .b(out_1285),
            .outp(out_1286)
        );        
        

        logic [WIDTH-1:0] out_1287;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1287 (
            .a(out_1285),
            .b(out_9),
            .outp(out_1287)
        );        
        

        logic [WIDTH-1:0] out_1288;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1288 (
            .a(out_1286),
            .b(out_1287),
            .outp(out_1288)
        );        
        

        logic [WIDTH-1:0] out_1289;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1289 (
            .a(out_1280),
            .b(out_1288),
            .outp(out_1289)
        );        
        

        logic [WIDTH-1:0] out_1290;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1290 (
            .a(out_1271),
            .b(out_1289),
            .outp(out_1290)
        );        
        

        logic [WIDTH-1:0] out_1291;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.35)
        ) inst_1291 (
            .outp(out_1291)
        );
        

        logic [WIDTH-1:0] out_1292;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1292 (
            .a(out_1291),
            .b(out_14),
            .outp(out_1292)
        );        
        

        logic [WIDTH-1:0] out_1293;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1293 (
            .a(out_1290),
            .b(out_1292),
            .outp(out_1293)
        );        
        

        logic [WIDTH-1:0] out_1294;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1294 (
            .a(out_1264),
            .b(out_1293),
            .outp(out_1294)
        );        
        

        logic [WIDTH-1:0] out_1295;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.523)
        ) inst_1295 (
            .outp(out_1295)
        );
        

        logic [WIDTH-1:0] out_1296;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1296 (
            .a(out_3),
            .b(out_1295),
            .outp(out_1296)
        );        
        

        logic [WIDTH-1:0] out_1297;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1297 (
            .in(out_1296),
            .outp(out_1297)
        );
        

        logic [WIDTH-1:0] out_1298;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.725)
        ) inst_1298 (
            .outp(out_1298)
        );
        

        logic [WIDTH-1:0] out_1299;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1299 (
            .a(out_1298),
            .b(out_14),
            .outp(out_1299)
        );        
        

        logic [WIDTH-1:0] out_1300;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1300 (
            .in(out_1299),
            .outp(out_1300)
        );
        

        logic [WIDTH-1:0] out_1301;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1301 (
            .a(out_1297),
            .b(out_1300),
            .outp(out_1301)
        );        
        

        logic [WIDTH-1:0] out_1302;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1302 (
            .in(out_1301),
            .outp(out_1302)
        );
        

        logic [WIDTH-1:0] out_1303;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1303 (
            .a(out_9),
            .b(out_1302),
            .outp(out_1303)
        );        
        

        logic [WIDTH-1:0] out_1304;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1304 (
            .a(out_1302),
            .b(out_21),
            .outp(out_1304)
        );        
        

        logic [WIDTH-1:0] out_1305;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1305 (
            .a(out_1303),
            .b(out_1304),
            .outp(out_1305)
        );        
        

        logic [WIDTH-1:0] out_1306;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1306 (
            .a(out_1294),
            .b(out_1305),
            .outp(out_1306)
        );        
        

        logic [WIDTH-1:0] out_1307;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0979996)
        ) inst_1307 (
            .outp(out_1307)
        );
        

        logic [WIDTH-1:0] out_1308;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1308 (
            .a(out_3),
            .b(out_1307),
            .outp(out_1308)
        );        
        

        logic [WIDTH-1:0] out_1309;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.00200015)
        ) inst_1309 (
            .outp(out_1309)
        );
        

        logic [WIDTH-1:0] out_1310;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1310 (
            .a(out_1309),
            .b(out_3),
            .outp(out_1310)
        );        
        

        logic [WIDTH-1:0] out_1311;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1311 (
            .in(out_1310),
            .outp(out_1311)
        );
        

        logic [WIDTH-1:0] out_1312;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1312 (
            .a(out_1308),
            .b(out_1311),
            .outp(out_1312)
        );        
        

        logic [WIDTH-1:0] out_1313;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1313 (
            .a(out_1312),
            .b(out_1244),
            .outp(out_1313)
        );        
        

        logic [WIDTH-1:0] out_1314;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1314 (
            .a(out_1313),
            .b(out_1299),
            .outp(out_1314)
        );        
        

        logic [WIDTH-1:0] out_1315;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1315 (
            .a(out_1306),
            .b(out_1314),
            .outp(out_1315)
        );        
        

        logic [WIDTH-1:0] out_1316;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.352)
        ) inst_1316 (
            .outp(out_1316)
        );
        

        logic [WIDTH-1:0] out_1317;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1317 (
            .a(out_1316),
            .b(out_3),
            .outp(out_1317)
        );        
        

        logic [WIDTH-1:0] out_1318;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.452)
        ) inst_1318 (
            .outp(out_1318)
        );
        

        logic [WIDTH-1:0] out_1319;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1319 (
            .a(out_1318),
            .b(out_3),
            .outp(out_1319)
        );        
        

        logic [WIDTH-1:0] out_1320;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1320 (
            .in(out_1319),
            .outp(out_1320)
        );
        

        logic [WIDTH-1:0] out_1321;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1321 (
            .a(out_1317),
            .b(out_1320),
            .outp(out_1321)
        );        
        

        logic [WIDTH-1:0] out_1322;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1322 (
            .a(out_1321),
            .b(out_1244),
            .outp(out_1322)
        );        
        

        logic [WIDTH-1:0] out_1323;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0)
        ) inst_1323 (
            .outp(out_1323)
        );
        

        logic [WIDTH-1:0] out_1324;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1324 (
            .a(out_1323),
            .b(out_14),
            .outp(out_1324)
        );        
        

        logic [WIDTH-1:0] out_1325;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1325 (
            .a(out_1322),
            .b(out_1324),
            .outp(out_1325)
        );        
        

        logic [WIDTH-1:0] out_1326;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1326 (
            .a(out_1315),
            .b(out_1325),
            .outp(out_1326)
        );        
        

        logic [WIDTH-1:0] out_1327;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1327 (
            .a(out_1308),
            .b(out_1320),
            .outp(out_1327)
        );        
        

        logic [WIDTH-1:0] out_1328;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.177)
        ) inst_1328 (
            .outp(out_1328)
        );
        

        logic [WIDTH-1:0] out_1329;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1329 (
            .a(out_1328),
            .b(out_3),
            .outp(out_1329)
        );        
        

        logic [WIDTH-1:0] out_1330;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1330 (
            .in(out_1329),
            .outp(out_1330)
        );
        

        logic [WIDTH-1:0] out_1331;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1331 (
            .a(out_1330),
            .b(out_1300),
            .outp(out_1331)
        );        
        

        logic [WIDTH-1:0] out_1332;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1332 (
            .in(out_1331),
            .outp(out_1332)
        );
        

        logic [WIDTH-1:0] out_1333;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1333 (
            .a(out_9),
            .b(out_1332),
            .outp(out_1333)
        );        
        

        logic [WIDTH-1:0] out_1334;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1334 (
            .a(out_1327),
            .b(out_1333),
            .outp(out_1334)
        );        
        

        logic [WIDTH-1:0] out_1335;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1335 (
            .a(out_1332),
            .b(out_21),
            .outp(out_1335)
        );        
        

        logic [WIDTH-1:0] out_1336;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1336 (
            .a(out_1334),
            .b(out_1335),
            .outp(out_1336)
        );        
        

        logic [WIDTH-1:0] out_1337;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.45)
        ) inst_1337 (
            .outp(out_1337)
        );
        

        logic [WIDTH-1:0] out_1338;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1338 (
            .a(out_1337),
            .b(out_14),
            .outp(out_1338)
        );        
        

        logic [WIDTH-1:0] out_1339;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1339 (
            .a(out_1336),
            .b(out_1338),
            .outp(out_1339)
        );        
        

        logic [WIDTH-1:0] out_1340;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.725)
        ) inst_1340 (
            .outp(out_1340)
        );
        

        logic [WIDTH-1:0] out_1341;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1341 (
            .a(out_1340),
            .b(out_14),
            .outp(out_1341)
        );        
        

        logic [WIDTH-1:0] out_1342;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1342 (
            .in(out_1341),
            .outp(out_1342)
        );
        

        logic [WIDTH-1:0] out_1343;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1343 (
            .a(out_1339),
            .b(out_1342),
            .outp(out_1343)
        );        
        

        logic [WIDTH-1:0] out_1344;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1344 (
            .a(out_1326),
            .b(out_1343),
            .outp(out_1344)
        );        
        

        logic [WIDTH-1:0] out_1345;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.4105)
        ) inst_1345 (
            .outp(out_1345)
        );
        

        logic [WIDTH-1:0] out_1346;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1346 (
            .a(out_3),
            .b(out_1345),
            .outp(out_1346)
        );        
        

        logic [WIDTH-1:0] out_1347;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1347 (
            .in(out_1346),
            .outp(out_1347)
        );
        

        logic [WIDTH-1:0] out_1348;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1348 (
            .a(out_1347),
            .b(out_1300),
            .outp(out_1348)
        );        
        

        logic [WIDTH-1:0] out_1349;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1349 (
            .in(out_1348),
            .outp(out_1349)
        );
        

        logic [WIDTH-1:0] out_1350;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1350 (
            .a(out_9),
            .b(out_1349),
            .outp(out_1350)
        );        
        

        logic [WIDTH-1:0] out_1351;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1351 (
            .a(out_1349),
            .b(out_21),
            .outp(out_1351)
        );        
        

        logic [WIDTH-1:0] out_1352;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1352 (
            .a(out_1350),
            .b(out_1351),
            .outp(out_1352)
        );        
        

        logic [WIDTH-1:0] out_1353;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1353 (
            .a(out_1352),
            .b(out_1338),
            .outp(out_1353)
        );        
        

        logic [WIDTH-1:0] out_1354;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6855)
        ) inst_1354 (
            .outp(out_1354)
        );
        

        logic [WIDTH-1:0] out_1355;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1355 (
            .a(out_3),
            .b(out_1354),
            .outp(out_1355)
        );        
        

        logic [WIDTH-1:0] out_1356;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1356 (
            .a(out_1353),
            .b(out_1355),
            .outp(out_1356)
        );        
        

        logic [WIDTH-1:0] out_1357;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1355)
        ) inst_1357 (
            .outp(out_1357)
        );
        

        logic [WIDTH-1:0] out_1358;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1358 (
            .a(out_1357),
            .b(out_3),
            .outp(out_1358)
        );        
        

        logic [WIDTH-1:0] out_1359;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1359 (
            .a(out_1356),
            .b(out_1358),
            .outp(out_1359)
        );        
        

        logic [WIDTH-1:0] out_1360;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.675)
        ) inst_1360 (
            .outp(out_1360)
        );
        

        logic [WIDTH-1:0] out_1361;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1361 (
            .a(out_1360),
            .b(out_14),
            .outp(out_1361)
        );        
        

        logic [WIDTH-1:0] out_1362;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1362 (
            .in(out_1361),
            .outp(out_1362)
        );
        

        logic [WIDTH-1:0] out_1363;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1363 (
            .a(out_1359),
            .b(out_1362),
            .outp(out_1363)
        );        
        

        logic [WIDTH-1:0] out_1364;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1364 (
            .a(out_1344),
            .b(out_1363),
            .outp(out_1364)
        );        
        

        logic [WIDTH-1:0] out_1365;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0105)
        ) inst_1365 (
            .outp(out_1365)
        );
        

        logic [WIDTH-1:0] out_1366;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1366 (
            .a(out_3),
            .b(out_1365),
            .outp(out_1366)
        );        
        

        logic [WIDTH-1:0] out_1367;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.9105)
        ) inst_1367 (
            .outp(out_1367)
        );
        

        logic [WIDTH-1:0] out_1368;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1368 (
            .a(out_1367),
            .b(out_3),
            .outp(out_1368)
        );        
        

        logic [WIDTH-1:0] out_1369;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1369 (
            .a(out_1366),
            .b(out_1368),
            .outp(out_1369)
        );        
        

        logic [WIDTH-1:0] out_1370;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1370 (
            .a(out_1369),
            .b(out_1244),
            .outp(out_1370)
        );        
        

        logic [WIDTH-1:0] out_1371;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1371 (
            .a(out_1370),
            .b(out_1338),
            .outp(out_1371)
        );        
        

        logic [WIDTH-1:0] out_1372;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1372 (
            .a(out_1364),
            .b(out_1371),
            .outp(out_1372)
        );        
        

        logic [WIDTH-1:0] out_1373;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.3)
        ) inst_1373 (
            .outp(out_1373)
        );
        

        logic [WIDTH-1:0] out_1374;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1374 (
            .a(out_1373),
            .b(out_14),
            .outp(out_1374)
        );        
        

        logic [WIDTH-1:0] out_1375;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1375 (
            .in(out_1374),
            .outp(out_1375)
        );
        

        logic [WIDTH-1:0] out_1376;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.9605)
        ) inst_1376 (
            .outp(out_1376)
        );
        

        logic [WIDTH-1:0] out_1377;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1377 (
            .a(out_3),
            .b(out_1376),
            .outp(out_1377)
        );        
        

        logic [WIDTH-1:0] out_1378;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1378 (
            .in(out_1377),
            .outp(out_1378)
        );
        

        logic [WIDTH-1:0] out_1379;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1379 (
            .a(out_1375),
            .b(out_1378),
            .outp(out_1379)
        );        
        

        logic [WIDTH-1:0] out_1380;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1380 (
            .in(out_1379),
            .outp(out_1380)
        );
        

        logic [WIDTH-1:0] out_1381;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1381 (
            .a(out_1380),
            .b(out_460),
            .outp(out_1381)
        );        
        

        logic [WIDTH-1:0] out_1382;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1382 (
            .a(out_1372),
            .b(out_1381),
            .outp(out_1382)
        );        
        

        logic [WIDTH-1:0] out_1383;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.775)
        ) inst_1383 (
            .outp(out_1383)
        );
        

        logic [WIDTH-1:0] out_1384;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1384 (
            .a(out_1383),
            .b(out_14),
            .outp(out_1384)
        );        
        

        logic [WIDTH-1:0] out_1385;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1385 (
            .in(out_1384),
            .outp(out_1385)
        );
        

        logic [WIDTH-1:0] out_1386;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6125)
        ) inst_1386 (
            .outp(out_1386)
        );
        

        logic [WIDTH-1:0] out_1387;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1387 (
            .a(out_1386),
            .b(out_14),
            .outp(out_1387)
        );        
        

        logic [WIDTH-1:0] out_1388;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1388 (
            .a(out_1385),
            .b(out_1387),
            .outp(out_1388)
        );        
        

        logic [WIDTH-1:0] out_1389;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.22783)
        ) inst_1389 (
            .outp(out_1389)
        );
        

        logic [WIDTH-1:0] out_1390;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1390 (
            .a(out_1389),
            .b(out_260),
            .outp(out_1390)
        );        
        

        logic [WIDTH-1:0] out_1391;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1391 (
            .a(out_1388),
            .b(out_1390),
            .outp(out_1391)
        );        
        

        logic [WIDTH-1:0] out_1392;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.39033)
        ) inst_1392 (
            .outp(out_1392)
        );
        

        logic [WIDTH-1:0] out_1393;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1393 (
            .a(out_260),
            .b(out_1392),
            .outp(out_1393)
        );        
        

        logic [WIDTH-1:0] out_1394;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1394 (
            .a(out_1391),
            .b(out_1393),
            .outp(out_1394)
        );        
        

        logic [WIDTH-1:0] out_1395;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.615)
        ) inst_1395 (
            .outp(out_1395)
        );
        

        logic [WIDTH-1:0] out_1396;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1396 (
            .a(out_1395),
            .b(out_14),
            .outp(out_1396)
        );        
        

        logic [WIDTH-1:0] out_1397;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1397 (
            .in(out_1396),
            .outp(out_1397)
        );
        

        logic [WIDTH-1:0] out_1398;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1398 (
            .in(out_1397),
            .outp(out_1398)
        );
        

        logic [WIDTH-1:0] out_1399;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.81689)
        ) inst_1399 (
            .outp(out_1399)
        );
        

        logic [WIDTH-1:0] out_1400;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1400 (
            .a(out_1399),
            .b(out_241),
            .outp(out_1400)
        );        
        

        logic [WIDTH-1:0] out_1401;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1401 (
            .in(out_1400),
            .outp(out_1401)
        );
        

        logic [WIDTH-1:0] out_1402;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1402 (
            .a(out_1398),
            .b(out_1401),
            .outp(out_1402)
        );        
        

        logic [WIDTH-1:0] out_1403;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1403 (
            .in(out_1402),
            .outp(out_1403)
        );
        

        logic [WIDTH-1:0] out_1404;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1404 (
            .a(out_1403),
            .b(out_250),
            .outp(out_1404)
        );        
        

        logic [WIDTH-1:0] out_1405;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1405 (
            .a(out_1394),
            .b(out_1404),
            .outp(out_1405)
        );        
        

        logic [WIDTH-1:0] out_1406;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1406 (
            .in(out_1405),
            .outp(out_1406)
        );
        

        logic [WIDTH-1:0] out_1407;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6125)
        ) inst_1407 (
            .outp(out_1407)
        );
        

        logic [WIDTH-1:0] out_1408;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1408 (
            .a(out_1407),
            .b(out_14),
            .outp(out_1408)
        );        
        

        logic [WIDTH-1:0] out_1409;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1409 (
            .in(out_1408),
            .outp(out_1409)
        );
        

        logic [WIDTH-1:0] out_1410;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1410 (
            .in(out_1409),
            .outp(out_1410)
        );
        

        logic [WIDTH-1:0] out_1411;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1411 (
            .in(out_1390),
            .outp(out_1411)
        );
        

        logic [WIDTH-1:0] out_1412;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1412 (
            .a(out_1410),
            .b(out_1411),
            .outp(out_1412)
        );        
        

        logic [WIDTH-1:0] out_1413;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1413 (
            .in(out_1412),
            .outp(out_1413)
        );
        

        logic [WIDTH-1:0] out_1414;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1414 (
            .a(out_1413),
            .b(out_275),
            .outp(out_1414)
        );        
        

        logic [WIDTH-1:0] out_1415;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1415 (
            .a(out_1406),
            .b(out_1414),
            .outp(out_1415)
        );        
        

        logic [WIDTH-1:0] out_1416;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1416 (
            .a(out_1382),
            .b(out_1415),
            .outp(out_1416)
        );        
        

        logic [WIDTH-1:0] out_1417;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8375)
        ) inst_1417 (
            .outp(out_1417)
        );
        

        logic [WIDTH-1:0] out_1418;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1418 (
            .a(out_1417),
            .b(out_14),
            .outp(out_1418)
        );        
        

        logic [WIDTH-1:0] out_1419;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1419 (
            .in(out_1418),
            .outp(out_1419)
        );
        

        logic [WIDTH-1:0] out_1420;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.22783)
        ) inst_1420 (
            .outp(out_1420)
        );
        

        logic [WIDTH-1:0] out_1421;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1421 (
            .a(out_260),
            .b(out_1420),
            .outp(out_1421)
        );        
        

        logic [WIDTH-1:0] out_1422;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1422 (
            .a(out_1419),
            .b(out_1421),
            .outp(out_1422)
        );        
        

        logic [WIDTH-1:0] out_1423;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.06533)
        ) inst_1423 (
            .outp(out_1423)
        );
        

        logic [WIDTH-1:0] out_1424;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1424 (
            .a(out_1423),
            .b(out_260),
            .outp(out_1424)
        );        
        

        logic [WIDTH-1:0] out_1425;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1425 (
            .a(out_1422),
            .b(out_1424),
            .outp(out_1425)
        );        
        

        logic [WIDTH-1:0] out_1426;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.675)
        ) inst_1426 (
            .outp(out_1426)
        );
        

        logic [WIDTH-1:0] out_1427;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1427 (
            .a(out_1426),
            .b(out_14),
            .outp(out_1427)
        );        
        

        logic [WIDTH-1:0] out_1428;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1428 (
            .a(out_1425),
            .b(out_1427),
            .outp(out_1428)
        );        
        

        logic [WIDTH-1:0] out_1429;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.835)
        ) inst_1429 (
            .outp(out_1429)
        );
        

        logic [WIDTH-1:0] out_1430;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1430 (
            .a(out_1429),
            .b(out_14),
            .outp(out_1430)
        );        
        

        logic [WIDTH-1:0] out_1431;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1431 (
            .in(out_1430),
            .outp(out_1431)
        );
        

        logic [WIDTH-1:0] out_1432;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.820223)
        ) inst_1432 (
            .outp(out_1432)
        );
        

        logic [WIDTH-1:0] out_1433;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1433 (
            .a(out_241),
            .b(out_1432),
            .outp(out_1433)
        );        
        

        logic [WIDTH-1:0] out_1434;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1434 (
            .in(out_1433),
            .outp(out_1434)
        );
        

        logic [WIDTH-1:0] out_1435;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1435 (
            .a(out_1431),
            .b(out_1434),
            .outp(out_1435)
        );        
        

        logic [WIDTH-1:0] out_1436;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1436 (
            .in(out_1435),
            .outp(out_1436)
        );
        

        logic [WIDTH-1:0] out_1437;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1437 (
            .a(out_1436),
            .b(out_250),
            .outp(out_1437)
        );        
        

        logic [WIDTH-1:0] out_1438;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1438 (
            .a(out_1428),
            .b(out_1437),
            .outp(out_1438)
        );        
        

        logic [WIDTH-1:0] out_1439;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1439 (
            .in(out_1438),
            .outp(out_1439)
        );
        

        logic [WIDTH-1:0] out_1440;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8375)
        ) inst_1440 (
            .outp(out_1440)
        );
        

        logic [WIDTH-1:0] out_1441;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1441 (
            .a(out_1440),
            .b(out_14),
            .outp(out_1441)
        );        
        

        logic [WIDTH-1:0] out_1442;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1442 (
            .in(out_1441),
            .outp(out_1442)
        );
        

        logic [WIDTH-1:0] out_1443;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1443 (
            .in(out_1421),
            .outp(out_1443)
        );
        

        logic [WIDTH-1:0] out_1444;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1444 (
            .a(out_1442),
            .b(out_1443),
            .outp(out_1444)
        );        
        

        logic [WIDTH-1:0] out_1445;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1445 (
            .in(out_1444),
            .outp(out_1445)
        );
        

        logic [WIDTH-1:0] out_1446;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1446 (
            .a(out_1445),
            .b(out_275),
            .outp(out_1446)
        );        
        

        logic [WIDTH-1:0] out_1447;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1447 (
            .a(out_1439),
            .b(out_1446),
            .outp(out_1447)
        );        
        

        logic [WIDTH-1:0] out_1448;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1448 (
            .a(out_1416),
            .b(out_1447),
            .outp(out_1448)
        );        
        

        logic [WIDTH-1:0] out_1449;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.207)
        ) inst_1449 (
            .outp(out_1449)
        );
        

        logic [WIDTH-1:0] out_1450;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1450 (
            .a(out_1449),
            .b(out_3),
            .outp(out_1450)
        );        
        

        logic [WIDTH-1:0] out_1451;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1451 (
            .in(out_1450),
            .outp(out_1451)
        );
        

        logic [WIDTH-1:0] out_1452;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1452 (
            .a(out_1451),
            .b(out_1300),
            .outp(out_1452)
        );        
        

        logic [WIDTH-1:0] out_1453;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1453 (
            .in(out_1452),
            .outp(out_1453)
        );
        

        logic [WIDTH-1:0] out_1454;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1454 (
            .a(out_9),
            .b(out_1453),
            .outp(out_1454)
        );        
        

        logic [WIDTH-1:0] out_1455;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1455 (
            .a(out_1453),
            .b(out_21),
            .outp(out_1455)
        );        
        

        logic [WIDTH-1:0] out_1456;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1456 (
            .a(out_1454),
            .b(out_1455),
            .outp(out_1456)
        );        
        

        logic [WIDTH-1:0] out_1457;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.932)
        ) inst_1457 (
            .outp(out_1457)
        );
        

        logic [WIDTH-1:0] out_1458;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1458 (
            .a(out_1457),
            .b(out_3),
            .outp(out_1458)
        );        
        

        logic [WIDTH-1:0] out_1459;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1459 (
            .a(out_1456),
            .b(out_1458),
            .outp(out_1459)
        );        
        

        logic [WIDTH-1:0] out_1460;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.482)
        ) inst_1460 (
            .outp(out_1460)
        );
        

        logic [WIDTH-1:0] out_1461;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1461 (
            .a(out_1460),
            .b(out_3),
            .outp(out_1461)
        );        
        

        logic [WIDTH-1:0] out_1462;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1462 (
            .in(out_1461),
            .outp(out_1462)
        );
        

        logic [WIDTH-1:0] out_1463;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1463 (
            .a(out_1459),
            .b(out_1462),
            .outp(out_1463)
        );        
        

        logic [WIDTH-1:0] out_1464;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1464 (
            .a(out_1463),
            .b(out_1338),
            .outp(out_1464)
        );        
        

        logic [WIDTH-1:0] out_1465;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1465 (
            .a(out_1464),
            .b(out_1362),
            .outp(out_1465)
        );        
        

        logic [WIDTH-1:0] out_1466;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1466 (
            .a(out_1448),
            .b(out_1465),
            .outp(out_1466)
        );        
        

        logic [WIDTH-1:0] out_1467;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.607)
        ) inst_1467 (
            .outp(out_1467)
        );
        

        logic [WIDTH-1:0] out_1468;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1468 (
            .a(out_1467),
            .b(out_3),
            .outp(out_1468)
        );        
        

        logic [WIDTH-1:0] out_1469;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.707)
        ) inst_1469 (
            .outp(out_1469)
        );
        

        logic [WIDTH-1:0] out_1470;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1470 (
            .a(out_1469),
            .b(out_3),
            .outp(out_1470)
        );        
        

        logic [WIDTH-1:0] out_1471;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1471 (
            .in(out_1470),
            .outp(out_1471)
        );
        

        logic [WIDTH-1:0] out_1472;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1472 (
            .a(out_1468),
            .b(out_1471),
            .outp(out_1472)
        );        
        

        logic [WIDTH-1:0] out_1473;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1473 (
            .a(out_1472),
            .b(out_1244),
            .outp(out_1473)
        );        
        

        logic [WIDTH-1:0] out_1474;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1474 (
            .a(out_1473),
            .b(out_1338),
            .outp(out_1474)
        );        
        

        logic [WIDTH-1:0] out_1475;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1475 (
            .a(out_1466),
            .b(out_1474),
            .outp(out_1475)
        );        
        

        logic [WIDTH-1:0] out_1476;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.657)
        ) inst_1476 (
            .outp(out_1476)
        );
        

        logic [WIDTH-1:0] out_1477;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1477 (
            .a(out_1476),
            .b(out_3),
            .outp(out_1477)
        );        
        

        logic [WIDTH-1:0] out_1478;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1478 (
            .in(out_1477),
            .outp(out_1478)
        );
        

        logic [WIDTH-1:0] out_1479;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1479 (
            .a(out_1375),
            .b(out_1478),
            .outp(out_1479)
        );        
        

        logic [WIDTH-1:0] out_1480;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1480 (
            .in(out_1479),
            .outp(out_1480)
        );
        

        logic [WIDTH-1:0] out_1481;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1481 (
            .a(out_1480),
            .b(out_460),
            .outp(out_1481)
        );        
        

        logic [WIDTH-1:0] out_1482;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1482 (
            .a(out_1475),
            .b(out_1481),
            .outp(out_1482)
        );        
        

        logic [WIDTH-1:0] out_1483;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.852)
        ) inst_1483 (
            .outp(out_1483)
        );
        

        logic [WIDTH-1:0] out_1484;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1484 (
            .a(out_1483),
            .b(out_3),
            .outp(out_1484)
        );        
        

        logic [WIDTH-1:0] out_1485;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1485 (
            .a(out_1235),
            .b(out_1484),
            .outp(out_1485)
        );        
        

        logic [WIDTH-1:0] out_1486;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.952)
        ) inst_1486 (
            .outp(out_1486)
        );
        

        logic [WIDTH-1:0] out_1487;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1487 (
            .a(out_1486),
            .b(out_3),
            .outp(out_1487)
        );        
        

        logic [WIDTH-1:0] out_1488;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1488 (
            .in(out_1487),
            .outp(out_1488)
        );
        

        logic [WIDTH-1:0] out_1489;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1489 (
            .a(out_1485),
            .b(out_1488),
            .outp(out_1489)
        );        
        

        logic [WIDTH-1:0] out_1490;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1490 (
            .a(out_1489),
            .b(out_1244),
            .outp(out_1490)
        );        
        

        logic [WIDTH-1:0] out_1491;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1491 (
            .a(out_1482),
            .b(out_1490),
            .outp(out_1491)
        );        
        

        logic [WIDTH-1:0] out_1492;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.35486)
        ) inst_1492 (
            .outp(out_1492)
        );
        

        logic [WIDTH-1:0] out_1493;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1493 (
            .a(out_1492),
            .b(out_3),
            .outp(out_1493)
        );        
        

        logic [WIDTH-1:0] out_1494;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.32288)
        ) inst_1494 (
            .outp(out_1494)
        );
        

        logic [WIDTH-1:0] out_1495;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1495 (
            .a(out_13),
            .b(out_1494),
            .outp(out_1495)
        );        
        

        logic [WIDTH-1:0] out_1496;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1496 (
            .a(out_1493),
            .b(out_1495),
            .outp(out_1496)
        );        
        

        logic [WIDTH-1:0] out_1497;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1497 (
            .in(out_1496),
            .outp(out_1497)
        );
        

        logic [WIDTH-1:0] out_1498;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1498 (
            .a(out_1497),
            .b(out_1300),
            .outp(out_1498)
        );        
        

        logic [WIDTH-1:0] out_1499;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1499 (
            .in(out_1498),
            .outp(out_1499)
        );
        

        logic [WIDTH-1:0] out_1500;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1500 (
            .a(out_9),
            .b(out_1499),
            .outp(out_1500)
        );        
        

        logic [WIDTH-1:0] out_1501;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1501 (
            .a(out_1499),
            .b(out_21),
            .outp(out_1501)
        );        
        

        logic [WIDTH-1:0] out_1502;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1502 (
            .a(out_1500),
            .b(out_1501),
            .outp(out_1502)
        );        
        

        logic [WIDTH-1:0] out_1503;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1503 (
            .a(out_1491),
            .b(out_1502),
            .outp(out_1503)
        );        
        

        logic [WIDTH-1:0] out_1504;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.662)
        ) inst_1504 (
            .outp(out_1504)
        );
        

        logic [WIDTH-1:0] out_1505;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1505 (
            .a(out_1504),
            .b(out_3),
            .outp(out_1505)
        );        
        

        logic [WIDTH-1:0] out_1506;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.762)
        ) inst_1506 (
            .outp(out_1506)
        );
        

        logic [WIDTH-1:0] out_1507;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1507 (
            .a(out_1506),
            .b(out_3),
            .outp(out_1507)
        );        
        

        logic [WIDTH-1:0] out_1508;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1508 (
            .in(out_1507),
            .outp(out_1508)
        );
        

        logic [WIDTH-1:0] out_1509;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1509 (
            .a(out_1505),
            .b(out_1508),
            .outp(out_1509)
        );        
        

        logic [WIDTH-1:0] out_1510;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1510 (
            .a(out_1509),
            .b(out_1324),
            .outp(out_1510)
        );        
        

        logic [WIDTH-1:0] out_1511;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.75)
        ) inst_1511 (
            .outp(out_1511)
        );
        

        logic [WIDTH-1:0] out_1512;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1512 (
            .a(out_1511),
            .b(out_14),
            .outp(out_1512)
        );        
        

        logic [WIDTH-1:0] out_1513;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1513 (
            .in(out_1512),
            .outp(out_1513)
        );
        

        logic [WIDTH-1:0] out_1514;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1514 (
            .a(out_1510),
            .b(out_1513),
            .outp(out_1514)
        );        
        

        logic [WIDTH-1:0] out_1515;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1515 (
            .a(out_1503),
            .b(out_1514),
            .outp(out_1515)
        );        
        

        logic [WIDTH-1:0] out_1516;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.512)
        ) inst_1516 (
            .outp(out_1516)
        );
        

        logic [WIDTH-1:0] out_1517;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1517 (
            .a(out_1516),
            .b(out_3),
            .outp(out_1517)
        );        
        

        logic [WIDTH-1:0] out_1518;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.912)
        ) inst_1518 (
            .outp(out_1518)
        );
        

        logic [WIDTH-1:0] out_1519;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1519 (
            .a(out_1518),
            .b(out_3),
            .outp(out_1519)
        );        
        

        logic [WIDTH-1:0] out_1520;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1520 (
            .in(out_1519),
            .outp(out_1520)
        );
        

        logic [WIDTH-1:0] out_1521;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1521 (
            .a(out_1517),
            .b(out_1520),
            .outp(out_1521)
        );        
        

        logic [WIDTH-1:0] out_1522;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1522 (
            .a(out_1521),
            .b(out_1292),
            .outp(out_1522)
        );        
        

        logic [WIDTH-1:0] out_1523;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.45)
        ) inst_1523 (
            .outp(out_1523)
        );
        

        logic [WIDTH-1:0] out_1524;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1524 (
            .a(out_1523),
            .b(out_14),
            .outp(out_1524)
        );        
        

        logic [WIDTH-1:0] out_1525;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1525 (
            .in(out_1524),
            .outp(out_1525)
        );
        

        logic [WIDTH-1:0] out_1526;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1526 (
            .a(out_1522),
            .b(out_1525),
            .outp(out_1526)
        );        
        

        logic [WIDTH-1:0] out_1527;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1527 (
            .a(out_1515),
            .b(out_1526),
            .outp(out_1527)
        );        
        

        logic [WIDTH-1:0] out_1528;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1528 (
            .in(out_1517),
            .outp(out_1528)
        );
        

        logic [WIDTH-1:0] out_1529;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1529 (
            .in(out_1512),
            .outp(out_1529)
        );
        

        logic [WIDTH-1:0] out_1530;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1530 (
            .a(out_1528),
            .b(out_1529),
            .outp(out_1530)
        );        
        

        logic [WIDTH-1:0] out_1531;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1531 (
            .in(out_1530),
            .outp(out_1531)
        );
        

        logic [WIDTH-1:0] out_1532;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1532 (
            .a(out_336),
            .b(out_1531),
            .outp(out_1532)
        );        
        

        logic [WIDTH-1:0] out_1533;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1533 (
            .a(out_1521),
            .b(out_1532),
            .outp(out_1533)
        );        
        

        logic [WIDTH-1:0] out_1534;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1534 (
            .a(out_1531),
            .b(out_343),
            .outp(out_1534)
        );        
        

        logic [WIDTH-1:0] out_1535;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1535 (
            .a(out_1533),
            .b(out_1534),
            .outp(out_1535)
        );        
        

        logic [WIDTH-1:0] out_1536;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1536 (
            .a(out_1535),
            .b(out_1244),
            .outp(out_1536)
        );        
        

        logic [WIDTH-1:0] out_1537;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1537 (
            .a(out_1536),
            .b(out_1512),
            .outp(out_1537)
        );        
        

        logic [WIDTH-1:0] out_1538;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1538 (
            .a(out_1527),
            .b(out_1537),
            .outp(out_1538)
        );        
        

        logic [WIDTH-1:0] out_1539;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.27)
        ) inst_1539 (
            .outp(out_1539)
        );
        

        logic [WIDTH-1:0] out_1540;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1540 (
            .a(out_1539),
            .b(out_3),
            .outp(out_1540)
        );        
        

        logic [WIDTH-1:0] out_1541;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.37)
        ) inst_1541 (
            .outp(out_1541)
        );
        

        logic [WIDTH-1:0] out_1542;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1542 (
            .a(out_1541),
            .b(out_3),
            .outp(out_1542)
        );        
        

        logic [WIDTH-1:0] out_1543;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1543 (
            .in(out_1542),
            .outp(out_1543)
        );
        

        logic [WIDTH-1:0] out_1544;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1544 (
            .a(out_1540),
            .b(out_1543),
            .outp(out_1544)
        );        
        

        logic [WIDTH-1:0] out_1545;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1545 (
            .a(out_1544),
            .b(out_1244),
            .outp(out_1545)
        );        
        

        logic [WIDTH-1:0] out_1546;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1546 (
            .a(out_1545),
            .b(out_1338),
            .outp(out_1546)
        );        
        

        logic [WIDTH-1:0] out_1547;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1547 (
            .a(out_1538),
            .b(out_1546),
            .outp(out_1547)
        );        
        

        logic [WIDTH-1:0] out_1548;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.702)
        ) inst_1548 (
            .outp(out_1548)
        );
        

        logic [WIDTH-1:0] out_1549;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1549 (
            .a(out_1548),
            .b(out_3),
            .outp(out_1549)
        );        
        

        logic [WIDTH-1:0] out_1550;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.802)
        ) inst_1550 (
            .outp(out_1550)
        );
        

        logic [WIDTH-1:0] out_1551;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1551 (
            .a(out_1550),
            .b(out_3),
            .outp(out_1551)
        );        
        

        logic [WIDTH-1:0] out_1552;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1552 (
            .in(out_1551),
            .outp(out_1552)
        );
        

        logic [WIDTH-1:0] out_1553;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1553 (
            .a(out_1549),
            .b(out_1552),
            .outp(out_1553)
        );        
        

        logic [WIDTH-1:0] out_1554;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1554 (
            .a(out_1553),
            .b(out_1324),
            .outp(out_1554)
        );        
        

        logic [WIDTH-1:0] out_1555;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1555 (
            .a(out_1554),
            .b(out_1513),
            .outp(out_1555)
        );        
        

        logic [WIDTH-1:0] out_1556;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1556 (
            .a(out_1547),
            .b(out_1555),
            .outp(out_1556)
        );        
        

        logic [WIDTH-1:0] out_1557;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.552)
        ) inst_1557 (
            .outp(out_1557)
        );
        

        logic [WIDTH-1:0] out_1558;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1558 (
            .a(out_1557),
            .b(out_3),
            .outp(out_1558)
        );        
        

        logic [WIDTH-1:0] out_1559;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.952)
        ) inst_1559 (
            .outp(out_1559)
        );
        

        logic [WIDTH-1:0] out_1560;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1560 (
            .a(out_1559),
            .b(out_3),
            .outp(out_1560)
        );        
        

        logic [WIDTH-1:0] out_1561;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1561 (
            .in(out_1560),
            .outp(out_1561)
        );
        

        logic [WIDTH-1:0] out_1562;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1562 (
            .a(out_1558),
            .b(out_1561),
            .outp(out_1562)
        );        
        

        logic [WIDTH-1:0] out_1563;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1563 (
            .a(out_1562),
            .b(out_1292),
            .outp(out_1563)
        );        
        

        logic [WIDTH-1:0] out_1564;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1564 (
            .a(out_1563),
            .b(out_1525),
            .outp(out_1564)
        );        
        

        logic [WIDTH-1:0] out_1565;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1565 (
            .a(out_1556),
            .b(out_1564),
            .outp(out_1565)
        );        
        

        logic [WIDTH-1:0] out_1566;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1566 (
            .in(out_1558),
            .outp(out_1566)
        );
        

        logic [WIDTH-1:0] out_1567;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1567 (
            .a(out_1566),
            .b(out_1529),
            .outp(out_1567)
        );        
        

        logic [WIDTH-1:0] out_1568;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1568 (
            .in(out_1567),
            .outp(out_1568)
        );
        

        logic [WIDTH-1:0] out_1569;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1569 (
            .a(out_336),
            .b(out_1568),
            .outp(out_1569)
        );        
        

        logic [WIDTH-1:0] out_1570;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1570 (
            .a(out_1562),
            .b(out_1569),
            .outp(out_1570)
        );        
        

        logic [WIDTH-1:0] out_1571;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1571 (
            .a(out_1568),
            .b(out_343),
            .outp(out_1571)
        );        
        

        logic [WIDTH-1:0] out_1572;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1572 (
            .a(out_1570),
            .b(out_1571),
            .outp(out_1572)
        );        
        

        logic [WIDTH-1:0] out_1573;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1573 (
            .a(out_1572),
            .b(out_1244),
            .outp(out_1573)
        );        
        

        logic [WIDTH-1:0] out_1574;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1574 (
            .a(out_1573),
            .b(out_1512),
            .outp(out_1574)
        );        
        

        logic [WIDTH-1:0] out_1575;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1575 (
            .a(out_1565),
            .b(out_1574),
            .outp(out_1575)
        );        
        

        logic [WIDTH-1:0] out_1576;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.072)
        ) inst_1576 (
            .outp(out_1576)
        );
        

        logic [WIDTH-1:0] out_1577;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1577 (
            .a(out_1576),
            .b(out_3),
            .outp(out_1577)
        );        
        

        logic [WIDTH-1:0] out_1578;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1578 (
            .a(out_1235),
            .b(out_1577),
            .outp(out_1578)
        );        
        

        logic [WIDTH-1:0] out_1579;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.172)
        ) inst_1579 (
            .outp(out_1579)
        );
        

        logic [WIDTH-1:0] out_1580;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1580 (
            .a(out_1579),
            .b(out_3),
            .outp(out_1580)
        );        
        

        logic [WIDTH-1:0] out_1581;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1581 (
            .in(out_1580),
            .outp(out_1581)
        );
        

        logic [WIDTH-1:0] out_1582;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1582 (
            .a(out_1578),
            .b(out_1581),
            .outp(out_1582)
        );        
        

        logic [WIDTH-1:0] out_1583;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1583 (
            .a(out_1582),
            .b(out_1244),
            .outp(out_1583)
        );        
        

        logic [WIDTH-1:0] out_1584;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1584 (
            .a(out_1575),
            .b(out_1583),
            .outp(out_1584)
        );        
        

        logic [WIDTH-1:0] out_1585;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.574857)
        ) inst_1585 (
            .outp(out_1585)
        );
        

        logic [WIDTH-1:0] out_1586;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1586 (
            .a(out_1585),
            .b(out_3),
            .outp(out_1586)
        );        
        

        logic [WIDTH-1:0] out_1587;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1587 (
            .a(out_1586),
            .b(out_1495),
            .outp(out_1587)
        );        
        

        logic [WIDTH-1:0] out_1588;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1588 (
            .in(out_1587),
            .outp(out_1588)
        );
        

        logic [WIDTH-1:0] out_1589;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1589 (
            .a(out_1588),
            .b(out_1300),
            .outp(out_1589)
        );        
        

        logic [WIDTH-1:0] out_1590;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1590 (
            .in(out_1589),
            .outp(out_1590)
        );
        

        logic [WIDTH-1:0] out_1591;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1591 (
            .a(out_9),
            .b(out_1590),
            .outp(out_1591)
        );        
        

        logic [WIDTH-1:0] out_1592;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1592 (
            .a(out_1590),
            .b(out_21),
            .outp(out_1592)
        );        
        

        logic [WIDTH-1:0] out_1593;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1593 (
            .a(out_1591),
            .b(out_1592),
            .outp(out_1593)
        );        
        

        logic [WIDTH-1:0] out_1594;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1594 (
            .a(out_1584),
            .b(out_1593),
            .outp(out_1594)
        );        
        

        logic [WIDTH-1:0] out_1595;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.25)
        ) inst_1595 (
            .outp(out_1595)
        );
        

        logic [WIDTH-1:0] out_1596;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1596 (
            .a(out_1595),
            .b(out_14),
            .outp(out_1596)
        );        
        

        logic [WIDTH-1:0] out_1597;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.882)
        ) inst_1597 (
            .outp(out_1597)
        );
        

        logic [WIDTH-1:0] out_1598;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1598 (
            .a(out_1597),
            .b(out_3),
            .outp(out_1598)
        );        
        

        logic [WIDTH-1:0] out_1599;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1599 (
            .a(out_1596),
            .b(out_1598),
            .outp(out_1599)
        );        
        

        logic [WIDTH-1:0] out_1600;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.982)
        ) inst_1600 (
            .outp(out_1600)
        );
        

        logic [WIDTH-1:0] out_1601;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1601 (
            .a(out_1600),
            .b(out_3),
            .outp(out_1601)
        );        
        

        logic [WIDTH-1:0] out_1602;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1602 (
            .in(out_1601),
            .outp(out_1602)
        );
        

        logic [WIDTH-1:0] out_1603;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1603 (
            .a(out_1599),
            .b(out_1602),
            .outp(out_1603)
        );        
        

        logic [WIDTH-1:0] out_1604;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1604 (
            .a(out_1603),
            .b(out_1244),
            .outp(out_1604)
        );        
        

        logic [WIDTH-1:0] out_1605;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1605 (
            .a(out_1594),
            .b(out_1604),
            .outp(out_1605)
        );        
        

        logic [WIDTH-1:0] out_1606;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.55)
        ) inst_1606 (
            .outp(out_1606)
        );
        

        logic [WIDTH-1:0] out_1607;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1607 (
            .a(out_1606),
            .b(out_14),
            .outp(out_1607)
        );        
        

        logic [WIDTH-1:0] out_1608;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1608 (
            .in(out_1607),
            .outp(out_1608)
        );
        

        logic [WIDTH-1:0] out_1609;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.732)
        ) inst_1609 (
            .outp(out_1609)
        );
        

        logic [WIDTH-1:0] out_1610;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1610 (
            .a(out_1609),
            .b(out_3),
            .outp(out_1610)
        );        
        

        logic [WIDTH-1:0] out_1611;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1611 (
            .a(out_1608),
            .b(out_1610),
            .outp(out_1611)
        );        
        

        logic [WIDTH-1:0] out_1612;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.132)
        ) inst_1612 (
            .outp(out_1612)
        );
        

        logic [WIDTH-1:0] out_1613;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1613 (
            .a(out_1612),
            .b(out_3),
            .outp(out_1613)
        );        
        

        logic [WIDTH-1:0] out_1614;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1614 (
            .in(out_1613),
            .outp(out_1614)
        );
        

        logic [WIDTH-1:0] out_1615;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1615 (
            .a(out_1611),
            .b(out_1614),
            .outp(out_1615)
        );        
        

        logic [WIDTH-1:0] out_1616;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1616 (
            .a(out_1615),
            .b(out_1338),
            .outp(out_1616)
        );        
        

        logic [WIDTH-1:0] out_1617;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1617 (
            .a(out_1605),
            .b(out_1616),
            .outp(out_1617)
        );        
        

        logic [WIDTH-1:0] out_1618;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1618 (
            .a(out_1610),
            .b(out_1614),
            .outp(out_1618)
        );        
        

        logic [WIDTH-1:0] out_1619;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1619 (
            .in(out_1596),
            .outp(out_1619)
        );
        

        logic [WIDTH-1:0] out_1620;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1620 (
            .a(out_1618),
            .b(out_1619),
            .outp(out_1620)
        );        
        

        logic [WIDTH-1:0] out_1621;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1621 (
            .in(out_1596),
            .outp(out_1621)
        );
        

        logic [WIDTH-1:0] out_1622;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1622 (
            .in(out_1610),
            .outp(out_1622)
        );
        

        logic [WIDTH-1:0] out_1623;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1623 (
            .a(out_1621),
            .b(out_1622),
            .outp(out_1623)
        );        
        

        logic [WIDTH-1:0] out_1624;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1624 (
            .in(out_1623),
            .outp(out_1624)
        );
        

        logic [WIDTH-1:0] out_1625;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1625 (
            .a(out_336),
            .b(out_1624),
            .outp(out_1625)
        );        
        

        logic [WIDTH-1:0] out_1626;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1626 (
            .a(out_1620),
            .b(out_1625),
            .outp(out_1626)
        );        
        

        logic [WIDTH-1:0] out_1627;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1627 (
            .a(out_1624),
            .b(out_343),
            .outp(out_1627)
        );        
        

        logic [WIDTH-1:0] out_1628;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1628 (
            .a(out_1626),
            .b(out_1627),
            .outp(out_1628)
        );        
        

        logic [WIDTH-1:0] out_1629;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1629 (
            .a(out_1628),
            .b(out_1324),
            .outp(out_1629)
        );        
        

        logic [WIDTH-1:0] out_1630;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1630 (
            .a(out_1617),
            .b(out_1629),
            .outp(out_1630)
        );        
        

        logic [WIDTH-1:0] out_1631;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.032)
        ) inst_1631 (
            .outp(out_1631)
        );
        

        logic [WIDTH-1:0] out_1632;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1632 (
            .a(out_1631),
            .b(out_3),
            .outp(out_1632)
        );        
        

        logic [WIDTH-1:0] out_1633;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1633 (
            .in(out_1632),
            .outp(out_1633)
        );
        

        logic [WIDTH-1:0] out_1634;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1634 (
            .a(out_1458),
            .b(out_1633),
            .outp(out_1634)
        );        
        

        logic [WIDTH-1:0] out_1635;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1635 (
            .a(out_1634),
            .b(out_1244),
            .outp(out_1635)
        );        
        

        logic [WIDTH-1:0] out_1636;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1636 (
            .a(out_1635),
            .b(out_1427),
            .outp(out_1636)
        );        
        

        logic [WIDTH-1:0] out_1637;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1637 (
            .a(out_1630),
            .b(out_1636),
            .outp(out_1637)
        );        
        

        logic [WIDTH-1:0] out_1638;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.382)
        ) inst_1638 (
            .outp(out_1638)
        );
        

        logic [WIDTH-1:0] out_1639;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1639 (
            .a(out_1638),
            .b(out_3),
            .outp(out_1639)
        );        
        

        logic [WIDTH-1:0] out_1640;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1640 (
            .a(out_1639),
            .b(out_1462),
            .outp(out_1640)
        );        
        

        logic [WIDTH-1:0] out_1641;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1641 (
            .a(out_1640),
            .b(out_1244),
            .outp(out_1641)
        );        
        

        logic [WIDTH-1:0] out_1642;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1642 (
            .a(out_1641),
            .b(out_1338),
            .outp(out_1642)
        );        
        

        logic [WIDTH-1:0] out_1643;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1643 (
            .a(out_1637),
            .b(out_1642),
            .outp(out_1643)
        );        
        

        logic [WIDTH-1:0] out_1644;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.25)
        ) inst_1644 (
            .outp(out_1644)
        );
        

        logic [WIDTH-1:0] out_1645;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1645 (
            .a(out_1644),
            .b(out_14),
            .outp(out_1645)
        );        
        

        logic [WIDTH-1:0] out_1646;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.35)
        ) inst_1646 (
            .outp(out_1646)
        );
        

        logic [WIDTH-1:0] out_1647;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1647 (
            .a(out_1646),
            .b(out_14),
            .outp(out_1647)
        );        
        

        logic [WIDTH-1:0] out_1648;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1648 (
            .in(out_1647),
            .outp(out_1648)
        );
        

        logic [WIDTH-1:0] out_1649;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1649 (
            .a(out_1645),
            .b(out_1648),
            .outp(out_1649)
        );        
        

        logic [WIDTH-1:0] out_1650;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.6385)
        ) inst_1650 (
            .outp(out_1650)
        );
        

        logic [WIDTH-1:0] out_1651;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1651 (
            .a(out_3),
            .b(out_1650),
            .outp(out_1651)
        );        
        

        logic [WIDTH-1:0] out_1652;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1652 (
            .a(out_1649),
            .b(out_1651),
            .outp(out_1652)
        );        
        

        logic [WIDTH-1:0] out_1653;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.2385)
        ) inst_1653 (
            .outp(out_1653)
        );
        

        logic [WIDTH-1:0] out_1654;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1654 (
            .a(out_1653),
            .b(out_3),
            .outp(out_1654)
        );        
        

        logic [WIDTH-1:0] out_1655;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1655 (
            .a(out_1652),
            .b(out_1654),
            .outp(out_1655)
        );        
        

        logic [WIDTH-1:0] out_1656;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1656 (
            .a(out_1643),
            .b(out_1655),
            .outp(out_1656)
        );        
        

        logic [WIDTH-1:0] out_1657;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1657 (
            .a(out_1651),
            .b(out_1654),
            .outp(out_1657)
        );        
        

        logic [WIDTH-1:0] out_1658;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.9)
        ) inst_1658 (
            .outp(out_1658)
        );
        

        logic [WIDTH-1:0] out_1659;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1659 (
            .a(out_1658),
            .b(out_14),
            .outp(out_1659)
        );        
        

        logic [WIDTH-1:0] out_1660;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1660 (
            .in(out_1659),
            .outp(out_1660)
        );
        

        logic [WIDTH-1:0] out_1661;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1661 (
            .a(out_1657),
            .b(out_1660),
            .outp(out_1661)
        );        
        

        logic [WIDTH-1:0] out_1662;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.65)
        ) inst_1662 (
            .outp(out_1662)
        );
        

        logic [WIDTH-1:0] out_1663;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1663 (
            .a(out_1662),
            .b(out_14),
            .outp(out_1663)
        );        
        

        logic [WIDTH-1:0] out_1664;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1664 (
            .in(out_1663),
            .outp(out_1664)
        );
        

        logic [WIDTH-1:0] out_1665;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1665 (
            .in(out_1651),
            .outp(out_1665)
        );
        

        logic [WIDTH-1:0] out_1666;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1666 (
            .a(out_1664),
            .b(out_1665),
            .outp(out_1666)
        );        
        

        logic [WIDTH-1:0] out_1667;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1667 (
            .in(out_1666),
            .outp(out_1667)
        );
        

        logic [WIDTH-1:0] out_1668;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1668 (
            .a(out_336),
            .b(out_1667),
            .outp(out_1668)
        );        
        

        logic [WIDTH-1:0] out_1669;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1669 (
            .a(out_1661),
            .b(out_1668),
            .outp(out_1669)
        );        
        

        logic [WIDTH-1:0] out_1670;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1670 (
            .a(out_1667),
            .b(out_343),
            .outp(out_1670)
        );        
        

        logic [WIDTH-1:0] out_1671;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1671 (
            .a(out_1669),
            .b(out_1670),
            .outp(out_1671)
        );        
        

        logic [WIDTH-1:0] out_1672;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1672 (
            .a(out_1671),
            .b(out_1663),
            .outp(out_1672)
        );        
        

        logic [WIDTH-1:0] out_1673;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1673 (
            .a(out_1656),
            .b(out_1672),
            .outp(out_1673)
        );        
        

        logic [WIDTH-1:0] out_1674;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.35)
        ) inst_1674 (
            .outp(out_1674)
        );
        

        logic [WIDTH-1:0] out_1675;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1675 (
            .a(out_1674),
            .b(out_14),
            .outp(out_1675)
        );        
        

        logic [WIDTH-1:0] out_1676;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1676 (
            .a(out_1660),
            .b(out_1675),
            .outp(out_1676)
        );        
        

        logic [WIDTH-1:0] out_1677;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.1135)
        ) inst_1677 (
            .outp(out_1677)
        );
        

        logic [WIDTH-1:0] out_1678;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1678 (
            .a(out_3),
            .b(out_1677),
            .outp(out_1678)
        );        
        

        logic [WIDTH-1:0] out_1679;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1679 (
            .a(out_1676),
            .b(out_1678),
            .outp(out_1679)
        );        
        

        logic [WIDTH-1:0] out_1680;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.0135)
        ) inst_1680 (
            .outp(out_1680)
        );
        

        logic [WIDTH-1:0] out_1681;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1681 (
            .a(out_1680),
            .b(out_3),
            .outp(out_1681)
        );        
        

        logic [WIDTH-1:0] out_1682;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1682 (
            .a(out_1679),
            .b(out_1681),
            .outp(out_1682)
        );        
        

        logic [WIDTH-1:0] out_1683;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1683 (
            .a(out_1673),
            .b(out_1682),
            .outp(out_1683)
        );        
        

        logic [WIDTH-1:0] out_1684;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2)
        ) inst_1684 (
            .outp(out_1684)
        );
        

        logic [WIDTH-1:0] out_1685;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1685 (
            .a(out_1684),
            .b(out_14),
            .outp(out_1685)
        );        
        

        logic [WIDTH-1:0] out_1686;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1686 (
            .in(out_1685),
            .outp(out_1686)
        );
        

        logic [WIDTH-1:0] out_1687;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.0635)
        ) inst_1687 (
            .outp(out_1687)
        );
        

        logic [WIDTH-1:0] out_1688;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1688 (
            .a(out_3),
            .b(out_1687),
            .outp(out_1688)
        );        
        

        logic [WIDTH-1:0] out_1689;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1689 (
            .in(out_1688),
            .outp(out_1689)
        );
        

        logic [WIDTH-1:0] out_1690;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1690 (
            .a(out_1686),
            .b(out_1689),
            .outp(out_1690)
        );        
        

        logic [WIDTH-1:0] out_1691;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1691 (
            .in(out_1690),
            .outp(out_1691)
        );
        

        logic [WIDTH-1:0] out_1692;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1692 (
            .a(out_1691),
            .b(out_460),
            .outp(out_1692)
        );        
        

        logic [WIDTH-1:0] out_1693;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1693 (
            .a(out_1683),
            .b(out_1692),
            .outp(out_1693)
        );        
        

        logic [WIDTH-1:0] out_1694;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.245)
        ) inst_1694 (
            .outp(out_1694)
        );
        

        logic [WIDTH-1:0] out_1695;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1695 (
            .a(out_1694),
            .b(out_152),
            .outp(out_1695)
        );        
        

        logic [WIDTH-1:0] out_1696;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1696 (
            .in(out_1695),
            .outp(out_1696)
        );
        

        logic [WIDTH-1:0] out_1697;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.15743)
        ) inst_1697 (
            .outp(out_1697)
        );
        

        logic [WIDTH-1:0] out_1698;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1698 (
            .a(out_1011),
            .b(out_1697),
            .outp(out_1698)
        );        
        

        logic [WIDTH-1:0] out_1699;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1699 (
            .a(out_127),
            .b(out_1698),
            .outp(out_1699)
        );        
        

        logic [WIDTH-1:0] out_1700;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1700 (
            .a(out_1696),
            .b(out_1699),
            .outp(out_1700)
        );        
        

        logic [WIDTH-1:0] out_1701;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.34743)
        ) inst_1701 (
            .outp(out_1701)
        );
        

        logic [WIDTH-1:0] out_1702;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1702 (
            .a(out_1017),
            .b(out_1701),
            .outp(out_1702)
        );        
        

        logic [WIDTH-1:0] out_1703;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1703 (
            .a(out_1702),
            .b(out_127),
            .outp(out_1703)
        );        
        

        logic [WIDTH-1:0] out_1704;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1704 (
            .a(out_1700),
            .b(out_1703),
            .outp(out_1704)
        );        
        

        logic [WIDTH-1:0] out_1705;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1705 (
            .a(out_1693),
            .b(out_1704),
            .outp(out_1705)
        );        
        

        logic [WIDTH-1:0] out_1706;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.34743)
        ) inst_1706 (
            .outp(out_1706)
        );
        

        logic [WIDTH-1:0] out_1707;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1707 (
            .a(out_1017),
            .b(out_1706),
            .outp(out_1707)
        );        
        

        logic [WIDTH-1:0] out_1708;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1708 (
            .a(out_127),
            .b(out_1707),
            .outp(out_1708)
        );        
        

        logic [WIDTH-1:0] out_1709;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1709 (
            .a(out_1695),
            .b(out_1708),
            .outp(out_1709)
        );        
        

        logic [WIDTH-1:0] out_1710;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1710 (
            .a(out_1698),
            .b(out_127),
            .outp(out_1710)
        );        
        

        logic [WIDTH-1:0] out_1711;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1711 (
            .a(out_1709),
            .b(out_1710),
            .outp(out_1711)
        );        
        

        logic [WIDTH-1:0] out_1712;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1712 (
            .a(out_1705),
            .b(out_1711),
            .outp(out_1712)
        );        
        

        logic [WIDTH-1:0] out_1713;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.19)
        ) inst_1713 (
            .outp(out_1713)
        );
        

        logic [WIDTH-1:0] out_1714;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1714 (
            .a(out_1713),
            .b(out_137),
            .outp(out_1714)
        );        
        

        logic [WIDTH-1:0] out_1715;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1715 (
            .a(out_1708),
            .b(out_1714),
            .outp(out_1715)
        );        
        

        logic [WIDTH-1:0] out_1716;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.10243)
        ) inst_1716 (
            .outp(out_1716)
        );
        

        logic [WIDTH-1:0] out_1717;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1717 (
            .a(out_1011),
            .b(out_1716),
            .outp(out_1717)
        );        
        

        logic [WIDTH-1:0] out_1718;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1718 (
            .a(out_1717),
            .b(out_127),
            .outp(out_1718)
        );        
        

        logic [WIDTH-1:0] out_1719;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1719 (
            .a(out_1715),
            .b(out_1718),
            .outp(out_1719)
        );        
        

        logic [WIDTH-1:0] out_1720;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1720 (
            .a(out_1712),
            .b(out_1719),
            .outp(out_1720)
        );        
        

        logic [WIDTH-1:0] out_1721;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1721 (
            .a(out_127),
            .b(out_1717),
            .outp(out_1721)
        );        
        

        logic [WIDTH-1:0] out_1722;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1722 (
            .a(out_1703),
            .b(out_1721),
            .outp(out_1722)
        );        
        

        logic [WIDTH-1:0] out_1723;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1723 (
            .in(out_1714),
            .outp(out_1723)
        );
        

        logic [WIDTH-1:0] out_1724;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1724 (
            .a(out_1722),
            .b(out_1723),
            .outp(out_1724)
        );        
        

        logic [WIDTH-1:0] out_1725;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1725 (
            .a(out_1720),
            .b(out_1724),
            .outp(out_1725)
        );        
        

        logic [WIDTH-1:0] out_1726;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1726 (
            .a(out_1713),
            .b(out_152),
            .outp(out_1726)
        );        
        

        logic [WIDTH-1:0] out_1727;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1727 (
            .in(out_1726),
            .outp(out_1727)
        );
        

        logic [WIDTH-1:0] out_1728;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1728 (
            .a(out_1699),
            .b(out_1727),
            .outp(out_1728)
        );        
        

        logic [WIDTH-1:0] out_1729;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.29243)
        ) inst_1729 (
            .outp(out_1729)
        );
        

        logic [WIDTH-1:0] out_1730;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1730 (
            .a(out_1017),
            .b(out_1729),
            .outp(out_1730)
        );        
        

        logic [WIDTH-1:0] out_1731;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1731 (
            .a(out_1730),
            .b(out_127),
            .outp(out_1731)
        );        
        

        logic [WIDTH-1:0] out_1732;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1732 (
            .a(out_1728),
            .b(out_1731),
            .outp(out_1732)
        );        
        

        logic [WIDTH-1:0] out_1733;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1733 (
            .a(out_1725),
            .b(out_1732),
            .outp(out_1733)
        );        
        

        logic [WIDTH-1:0] out_1734;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1734 (
            .a(out_1710),
            .b(out_1726),
            .outp(out_1734)
        );        
        

        logic [WIDTH-1:0] out_1735;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1735 (
            .a(out_127),
            .b(out_1730),
            .outp(out_1735)
        );        
        

        logic [WIDTH-1:0] out_1736;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1736 (
            .a(out_1734),
            .b(out_1735),
            .outp(out_1736)
        );        
        

        logic [WIDTH-1:0] out_1737;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1737 (
            .a(out_1733),
            .b(out_1736),
            .outp(out_1737)
        );        
        

        logic [WIDTH-1:0] out_1738;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1738 (
            .a(out_1718),
            .b(out_1735),
            .outp(out_1738)
        );        
        

        logic [WIDTH-1:0] out_1739;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.135)
        ) inst_1739 (
            .outp(out_1739)
        );
        

        logic [WIDTH-1:0] out_1740;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1740 (
            .a(out_1739),
            .b(out_137),
            .outp(out_1740)
        );        
        

        logic [WIDTH-1:0] out_1741;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1741 (
            .a(out_1738),
            .b(out_1740),
            .outp(out_1741)
        );        
        

        logic [WIDTH-1:0] out_1742;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1742 (
            .a(out_1737),
            .b(out_1741),
            .outp(out_1742)
        );        
        

        logic [WIDTH-1:0] out_1743;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1743 (
            .a(out_1721),
            .b(out_1731),
            .outp(out_1743)
        );        
        

        logic [WIDTH-1:0] out_1744;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1744 (
            .in(out_1740),
            .outp(out_1744)
        );
        

        logic [WIDTH-1:0] out_1745;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1745 (
            .a(out_1743),
            .b(out_1744),
            .outp(out_1745)
        );        
        

        logic [WIDTH-1:0] out_1746;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1746 (
            .a(out_1742),
            .b(out_1745),
            .outp(out_1746)
        );        
        

        logic [WIDTH-1:0] out_1747;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.24743)
        ) inst_1747 (
            .outp(out_1747)
        );
        

        logic [WIDTH-1:0] out_1748;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1748 (
            .a(out_1011),
            .b(out_127),
            .outp(out_1748)
        );        
        

        logic [WIDTH-1:0] out_1749;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1749 (
            .a(out_1747),
            .b(out_1748),
            .outp(out_1749)
        );        
        

        logic [WIDTH-1:0] out_1750;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1750 (
            .a(out_1727),
            .b(out_1749),
            .outp(out_1750)
        );        
        

        logic [WIDTH-1:0] out_1751;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1751 (
            .a(out_1017),
            .b(out_127),
            .outp(out_1751)
        );        
        

        logic [WIDTH-1:0] out_1752;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.11243)
        ) inst_1752 (
            .outp(out_1752)
        );
        

        logic [WIDTH-1:0] out_1753;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1753 (
            .a(out_1751),
            .b(out_1752),
            .outp(out_1753)
        );        
        

        logic [WIDTH-1:0] out_1754;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1754 (
            .a(out_1750),
            .b(out_1753),
            .outp(out_1754)
        );        
        

        logic [WIDTH-1:0] out_1755;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1755 (
            .a(out_1746),
            .b(out_1754),
            .outp(out_1755)
        );        
        

        logic [WIDTH-1:0] out_1756;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.12143)
        ) inst_1756 (
            .outp(out_1756)
        );
        

        logic [WIDTH-1:0] out_1757;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1757 (
            .a(out_1756),
            .b(out_194),
            .outp(out_1757)
        );        
        

        logic [WIDTH-1:0] out_1758;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.67143)
        ) inst_1758 (
            .outp(out_1758)
        );
        

        logic [WIDTH-1:0] out_1759;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1759 (
            .a(out_1758),
            .b(out_194),
            .outp(out_1759)
        );        
        

        logic [WIDTH-1:0] out_1760;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1760 (
            .in(out_1759),
            .outp(out_1760)
        );
        

        logic [WIDTH-1:0] out_1761;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1761 (
            .a(out_1757),
            .b(out_1760),
            .outp(out_1761)
        );        
        

        logic [WIDTH-1:0] out_1762;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1762 (
            .in(out_1243),
            .outp(out_1762)
        );
        

        logic [WIDTH-1:0] out_1763;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.90179)
        ) inst_1763 (
            .outp(out_1763)
        );
        

        logic [WIDTH-1:0] out_1764;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1764 (
            .a(out_1763),
            .b(out_204),
            .outp(out_1764)
        );        
        

        logic [WIDTH-1:0] out_1765;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1765 (
            .in(out_1764),
            .outp(out_1765)
        );
        

        logic [WIDTH-1:0] out_1766;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1766 (
            .a(out_1762),
            .b(out_1765),
            .outp(out_1766)
        );        
        

        logic [WIDTH-1:0] out_1767;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1767 (
            .in(out_1766),
            .outp(out_1767)
        );
        

        logic [WIDTH-1:0] out_1768;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1768 (
            .a(out_200),
            .b(out_1767),
            .outp(out_1768)
        );        
        

        logic [WIDTH-1:0] out_1769;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1769 (
            .a(out_1761),
            .b(out_1768),
            .outp(out_1769)
        );        
        

        logic [WIDTH-1:0] out_1770;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1770 (
            .in(out_1757),
            .outp(out_1770)
        );
        

        logic [WIDTH-1:0] out_1771;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1771 (
            .a(out_1762),
            .b(out_1770),
            .outp(out_1771)
        );        
        

        logic [WIDTH-1:0] out_1772;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1772 (
            .in(out_1771),
            .outp(out_1772)
        );
        

        logic [WIDTH-1:0] out_1773;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1773 (
            .a(out_1772),
            .b(out_214),
            .outp(out_1773)
        );        
        

        logic [WIDTH-1:0] out_1774;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1774 (
            .a(out_1769),
            .b(out_1773),
            .outp(out_1774)
        );        
        

        logic [WIDTH-1:0] out_1775;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1775 (
            .a(out_1774),
            .b(out_1244),
            .outp(out_1775)
        );        
        

        logic [WIDTH-1:0] out_1776;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1776 (
            .a(out_1775),
            .b(out_1338),
            .outp(out_1776)
        );        
        

        logic [WIDTH-1:0] out_1777;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1777 (
            .a(out_1755),
            .b(out_1776),
            .outp(out_1777)
        );        
        

        logic [WIDTH-1:0] out_1778;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.47)
        ) inst_1778 (
            .outp(out_1778)
        );
        

        logic [WIDTH-1:0] out_1779;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1779 (
            .a(out_1778),
            .b(out_3),
            .outp(out_1779)
        );        
        

        logic [WIDTH-1:0] out_1780;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.97)
        ) inst_1780 (
            .outp(out_1780)
        );
        

        logic [WIDTH-1:0] out_1781;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1781 (
            .a(out_1780),
            .b(out_3),
            .outp(out_1781)
        );        
        

        logic [WIDTH-1:0] out_1782;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1782 (
            .in(out_1781),
            .outp(out_1782)
        );
        

        logic [WIDTH-1:0] out_1783;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1783 (
            .a(out_1779),
            .b(out_1782),
            .outp(out_1783)
        );        
        

        logic [WIDTH-1:0] out_1784;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.685)
        ) inst_1784 (
            .outp(out_1784)
        );
        

        logic [WIDTH-1:0] out_1785;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1785 (
            .a(out_1784),
            .b(out_14),
            .outp(out_1785)
        );        
        

        logic [WIDTH-1:0] out_1786;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1786 (
            .a(out_1783),
            .b(out_1785),
            .outp(out_1786)
        );        
        

        logic [WIDTH-1:0] out_1787;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.775)
        ) inst_1787 (
            .outp(out_1787)
        );
        

        logic [WIDTH-1:0] out_1788;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1788 (
            .a(out_1787),
            .b(out_14),
            .outp(out_1788)
        );        
        

        logic [WIDTH-1:0] out_1789;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1789 (
            .in(out_1788),
            .outp(out_1789)
        );
        

        logic [WIDTH-1:0] out_1790;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1790 (
            .a(out_1786),
            .b(out_1789),
            .outp(out_1790)
        );        
        

        logic [WIDTH-1:0] out_1791;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.745)
        ) inst_1791 (
            .outp(out_1791)
        );
        

        logic [WIDTH-1:0] out_1792;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1792 (
            .a(out_1791),
            .b(out_3),
            .outp(out_1792)
        );        
        

        logic [WIDTH-1:0] out_1793;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1793 (
            .in(out_1792),
            .outp(out_1793)
        );
        

        logic [WIDTH-1:0] out_1794;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1794 (
            .a(out_1793),
            .b(out_1300),
            .outp(out_1794)
        );        
        

        logic [WIDTH-1:0] out_1795;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1795 (
            .in(out_1794),
            .outp(out_1795)
        );
        

        logic [WIDTH-1:0] out_1796;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1796 (
            .a(out_1795),
            .b(out_21),
            .outp(out_1796)
        );        
        

        logic [WIDTH-1:0] out_1797;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.0405)
        ) inst_1797 (
            .outp(out_1797)
        );
        

        logic [WIDTH-1:0] out_1798;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1798 (
            .a(out_1797),
            .b(out_556),
            .outp(out_1798)
        );        
        

        logic [WIDTH-1:0] out_1799;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1799 (
            .a(out_1798),
            .b(out_559),
            .outp(out_1799)
        );        
        

        logic [WIDTH-1:0] out_1800;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.9905)
        ) inst_1800 (
            .outp(out_1800)
        );
        

        logic [WIDTH-1:0] out_1801;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1801 (
            .a(out_556),
            .b(out_1800),
            .outp(out_1801)
        );        
        

        logic [WIDTH-1:0] out_1802;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1802 (
            .a(out_1801),
            .b(out_566),
            .outp(out_1802)
        );        
        

        logic [WIDTH-1:0] out_1803;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1803 (
            .in(out_1802),
            .outp(out_1803)
        );
        

        logic [WIDTH-1:0] out_1804;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1804 (
            .a(out_1799),
            .b(out_1803),
            .outp(out_1804)
        );        
        

        logic [WIDTH-1:0] out_1805;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.77125)
        ) inst_1805 (
            .outp(out_1805)
        );
        

        logic [WIDTH-1:0] out_1806;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1806 (
            .a(out_1805),
            .b(out_553),
            .outp(out_1806)
        );        
        

        logic [WIDTH-1:0] out_1807;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1807 (
            .a(out_1804),
            .b(out_1806),
            .outp(out_1807)
        );        
        

        logic [WIDTH-1:0] out_1808;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.9905)
        ) inst_1808 (
            .outp(out_1808)
        );
        

        logic [WIDTH-1:0] out_1809;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1809 (
            .a(out_556),
            .b(out_1808),
            .outp(out_1809)
        );        
        

        logic [WIDTH-1:0] out_1810;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1810 (
            .a(out_1809),
            .b(out_566),
            .outp(out_1810)
        );        
        

        logic [WIDTH-1:0] out_1811;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1811 (
            .a(out_559),
            .b(out_1798),
            .outp(out_1811)
        );        
        

        logic [WIDTH-1:0] out_1812;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1812 (
            .a(out_1810),
            .b(out_1811),
            .outp(out_1812)
        );        
        

        logic [WIDTH-1:0] out_1813;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1813 (
            .in(out_1806),
            .outp(out_1813)
        );
        

        logic [WIDTH-1:0] out_1814;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1814 (
            .a(out_1812),
            .b(out_1813),
            .outp(out_1814)
        );        
        

        logic [WIDTH-1:0] out_1815;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1815 (
            .a(out_1807),
            .b(out_1814),
            .outp(out_1815)
        );        
        

        logic [WIDTH-1:0] out_1816;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1816 (
            .in(out_1815),
            .outp(out_1816)
        );
        

        logic [WIDTH-1:0] out_1817;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1817 (
            .a(out_1796),
            .b(out_1816),
            .outp(out_1817)
        );        
        

        logic [WIDTH-1:0] out_1818;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1818 (
            .a(out_9),
            .b(out_1795),
            .outp(out_1818)
        );        
        

        logic [WIDTH-1:0] out_1819;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1819 (
            .a(out_1817),
            .b(out_1818),
            .outp(out_1819)
        );        
        

        logic [WIDTH-1:0] out_1820;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1820 (
            .a(out_1790),
            .b(out_1819),
            .outp(out_1820)
        );        
        

        logic [WIDTH-1:0] out_1821;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1821 (
            .a(out_1796),
            .b(out_1820),
            .outp(out_1821)
        );        
        

        logic [WIDTH-1:0] out_1822;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1822 (
            .a(out_1777),
            .b(out_1821),
            .outp(out_1822)
        );        
        

        logic [WIDTH-1:0] out_1823;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1823 (
            .a(out_13),
            .b(out_555),
            .outp(out_1823)
        );        
        

        logic [WIDTH-1:0] out_1824;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.02163)
        ) inst_1824 (
            .outp(out_1824)
        );
        

        logic [WIDTH-1:0] out_1825;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.27642)
        ) inst_1825 (
            .outp(out_1825)
        );
        

        logic [WIDTH-1:0] out_1826;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1826 (
            .a(out_1),
            .b(out_1825),
            .outp(out_1826)
        );        
        

        logic [WIDTH-1:0] out_1827;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1827 (
            .a(out_1824),
            .b(out_1826),
            .outp(out_1827)
        );        
        

        logic [WIDTH-1:0] out_1828;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1828 (
            .a(out_1823),
            .b(out_1827),
            .outp(out_1828)
        );        
        

        logic [WIDTH-1:0] out_1829;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.35775)
        ) inst_1829 (
            .outp(out_1829)
        );
        

        logic [WIDTH-1:0] out_1830;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5122)
        ) inst_1830 (
            .outp(out_1830)
        );
        

        logic [WIDTH-1:0] out_1831;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1831 (
            .a(out_1),
            .b(out_1830),
            .outp(out_1831)
        );        
        

        logic [WIDTH-1:0] out_1832;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1832 (
            .a(out_1829),
            .b(out_1831),
            .outp(out_1832)
        );        
        

        logic [WIDTH-1:0] out_1833;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1833 (
            .a(out_1828),
            .b(out_1832),
            .outp(out_1833)
        );        
        

        logic [WIDTH-1:0] out_1834;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1834 (
            .a(out_867),
            .b(out_555),
            .outp(out_1834)
        );        
        

        logic [WIDTH-1:0] out_1835;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.48875)
        ) inst_1835 (
            .outp(out_1835)
        );
        

        logic [WIDTH-1:0] out_1836;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1836 (
            .a(out_1834),
            .b(out_1835),
            .outp(out_1836)
        );        
        

        logic [WIDTH-1:0] out_1837;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1837 (
            .in(out_1836),
            .outp(out_1837)
        );
        

        logic [WIDTH-1:0] out_1838;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1838 (
            .a(out_1833),
            .b(out_1837),
            .outp(out_1838)
        );        
        

        logic [WIDTH-1:0] out_1839;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.48875)
        ) inst_1839 (
            .outp(out_1839)
        );
        

        logic [WIDTH-1:0] out_1840;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1840 (
            .a(out_1834),
            .b(out_1839),
            .outp(out_1840)
        );        
        

        logic [WIDTH-1:0] out_1841;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1841 (
            .in(out_1832),
            .outp(out_1841)
        );
        

        logic [WIDTH-1:0] out_1842;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1842 (
            .a(out_1840),
            .b(out_1841),
            .outp(out_1842)
        );        
        

        logic [WIDTH-1:0] out_1843;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.02162)
        ) inst_1843 (
            .outp(out_1843)
        );
        

        logic [WIDTH-1:0] out_1844;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1844 (
            .a(out_1843),
            .b(out_1826),
            .outp(out_1844)
        );        
        

        logic [WIDTH-1:0] out_1845;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1845 (
            .a(out_1844),
            .b(out_1823),
            .outp(out_1845)
        );        
        

        logic [WIDTH-1:0] out_1846;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1846 (
            .a(out_1842),
            .b(out_1845),
            .outp(out_1846)
        );        
        

        logic [WIDTH-1:0] out_1847;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1847 (
            .a(out_1838),
            .b(out_1846),
            .outp(out_1847)
        );        
        

        logic [WIDTH-1:0] out_1848;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1848 (
            .in(out_1847),
            .outp(out_1848)
        );
        

        logic [WIDTH-1:0] out_1849;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.325)
        ) inst_1849 (
            .outp(out_1849)
        );
        

        logic [WIDTH-1:0] out_1850;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1850 (
            .a(out_1849),
            .b(out_3),
            .outp(out_1850)
        );        
        

        logic [WIDTH-1:0] out_1851;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1851 (
            .in(out_1850),
            .outp(out_1851)
        );
        

        logic [WIDTH-1:0] out_1852;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1852 (
            .a(out_1851),
            .b(out_1300),
            .outp(out_1852)
        );        
        

        logic [WIDTH-1:0] out_1853;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1853 (
            .in(out_1852),
            .outp(out_1853)
        );
        

        logic [WIDTH-1:0] out_1854;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1854 (
            .a(out_9),
            .b(out_1853),
            .outp(out_1854)
        );        
        

        logic [WIDTH-1:0] out_1855;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1855 (
            .a(out_1848),
            .b(out_1854),
            .outp(out_1855)
        );        
        

        logic [WIDTH-1:0] out_1856;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1856 (
            .a(out_1853),
            .b(out_21),
            .outp(out_1856)
        );        
        

        logic [WIDTH-1:0] out_1857;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1857 (
            .a(out_1855),
            .b(out_1856),
            .outp(out_1857)
        );        
        

        logic [WIDTH-1:0] out_1858;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1858 (
            .a(out_1822),
            .b(out_1857),
            .outp(out_1858)
        );        
        

        logic [WIDTH-1:0] out_1859;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.9)
        ) inst_1859 (
            .outp(out_1859)
        );
        

        logic [WIDTH-1:0] out_1860;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1860 (
            .a(out_1859),
            .b(out_14),
            .outp(out_1860)
        );        
        

        logic [WIDTH-1:0] out_1861;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1861 (
            .in(out_1663),
            .outp(out_1861)
        );
        

        logic [WIDTH-1:0] out_1862;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1862 (
            .a(out_1860),
            .b(out_1861),
            .outp(out_1862)
        );        
        

        logic [WIDTH-1:0] out_1863;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.4885)
        ) inst_1863 (
            .outp(out_1863)
        );
        

        logic [WIDTH-1:0] out_1864;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1864 (
            .a(out_3),
            .b(out_1863),
            .outp(out_1864)
        );        
        

        logic [WIDTH-1:0] out_1865;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1865 (
            .a(out_1862),
            .b(out_1864),
            .outp(out_1865)
        );        
        

        logic [WIDTH-1:0] out_1866;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.3885)
        ) inst_1866 (
            .outp(out_1866)
        );
        

        logic [WIDTH-1:0] out_1867;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1867 (
            .a(out_1866),
            .b(out_3),
            .outp(out_1867)
        );        
        

        logic [WIDTH-1:0] out_1868;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1868 (
            .a(out_1865),
            .b(out_1867),
            .outp(out_1868)
        );        
        

        logic [WIDTH-1:0] out_1869;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1869 (
            .a(out_1858),
            .b(out_1868),
            .outp(out_1869)
        );        
        

        logic [WIDTH-1:0] out_1870;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1870 (
            .a(out_1660),
            .b(out_1860),
            .outp(out_1870)
        );        
        

        logic [WIDTH-1:0] out_1871;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.625)
        ) inst_1871 (
            .outp(out_1871)
        );
        

        logic [WIDTH-1:0] out_1872;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1872 (
            .a(out_1871),
            .b(out_14),
            .outp(out_1872)
        );        
        

        logic [WIDTH-1:0] out_1873;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1873 (
            .in(out_1872),
            .outp(out_1873)
        );
        

        logic [WIDTH-1:0] out_1874;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1805)
        ) inst_1874 (
            .outp(out_1874)
        );
        

        logic [WIDTH-1:0] out_1875;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1875 (
            .a(out_3),
            .b(out_1874),
            .outp(out_1875)
        );        
        

        logic [WIDTH-1:0] out_1876;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1876 (
            .in(out_1875),
            .outp(out_1876)
        );
        

        logic [WIDTH-1:0] out_1877;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1877 (
            .a(out_1873),
            .b(out_1876),
            .outp(out_1877)
        );        
        

        logic [WIDTH-1:0] out_1878;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1878 (
            .in(out_1877),
            .outp(out_1878)
        );
        

        logic [WIDTH-1:0] out_1879;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1879 (
            .a(out_9),
            .b(out_1878),
            .outp(out_1879)
        );        
        

        logic [WIDTH-1:0] out_1880;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1880 (
            .a(out_1870),
            .b(out_1879),
            .outp(out_1880)
        );        
        

        logic [WIDTH-1:0] out_1881;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1881 (
            .a(out_1878),
            .b(out_21),
            .outp(out_1881)
        );        
        

        logic [WIDTH-1:0] out_1882;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1882 (
            .a(out_1880),
            .b(out_1881),
            .outp(out_1882)
        );        
        

        logic [WIDTH-1:0] out_1883;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.9055)
        ) inst_1883 (
            .outp(out_1883)
        );
        

        logic [WIDTH-1:0] out_1884;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1884 (
            .a(out_3),
            .b(out_1883),
            .outp(out_1884)
        );        
        

        logic [WIDTH-1:0] out_1885;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1885 (
            .a(out_1882),
            .b(out_1884),
            .outp(out_1885)
        );        
        

        logic [WIDTH-1:0] out_1886;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1805)
        ) inst_1886 (
            .outp(out_1886)
        );
        

        logic [WIDTH-1:0] out_1887;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1887 (
            .a(out_1886),
            .b(out_3),
            .outp(out_1887)
        );        
        

        logic [WIDTH-1:0] out_1888;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1888 (
            .a(out_1885),
            .b(out_1887),
            .outp(out_1888)
        );        
        

        logic [WIDTH-1:0] out_1889;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1889 (
            .a(out_1869),
            .b(out_1888),
            .outp(out_1889)
        );        
        

        logic [WIDTH-1:0] out_1890;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.84553)
        ) inst_1890 (
            .outp(out_1890)
        );
        

        logic [WIDTH-1:0] out_1891;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1891 (
            .a(out_1),
            .b(out_1890),
            .outp(out_1891)
        );        
        

        logic [WIDTH-1:0] out_1892;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.880675)
        ) inst_1892 (
            .outp(out_1892)
        );
        

        logic [WIDTH-1:0] out_1893;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1893 (
            .a(out_137),
            .b(out_1892),
            .outp(out_1893)
        );        
        

        logic [WIDTH-1:0] out_1894;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1894 (
            .a(out_1891),
            .b(out_1893),
            .outp(out_1894)
        );        
        

        logic [WIDTH-1:0] out_1895;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.590637)
        ) inst_1895 (
            .outp(out_1895)
        );
        

        logic [WIDTH-1:0] out_1896;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.82927)
        ) inst_1896 (
            .outp(out_1896)
        );
        

        logic [WIDTH-1:0] out_1897;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1897 (
            .a(out_1),
            .b(out_1896),
            .outp(out_1897)
        );        
        

        logic [WIDTH-1:0] out_1898;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1898 (
            .a(out_1895),
            .b(out_1897),
            .outp(out_1898)
        );        
        

        logic [WIDTH-1:0] out_1899;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1899 (
            .a(out_1898),
            .b(out_566),
            .outp(out_1899)
        );        
        

        logic [WIDTH-1:0] out_1900;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1900 (
            .in(out_1899),
            .outp(out_1900)
        );
        

        logic [WIDTH-1:0] out_1901;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1901 (
            .a(out_1894),
            .b(out_1900),
            .outp(out_1901)
        );        
        

        logic [WIDTH-1:0] out_1902;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.27381)
        ) inst_1902 (
            .outp(out_1902)
        );
        

        logic [WIDTH-1:0] out_1903;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.87805)
        ) inst_1903 (
            .outp(out_1903)
        );
        

        logic [WIDTH-1:0] out_1904;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1904 (
            .a(out_13),
            .b(out_1903),
            .outp(out_1904)
        );        
        

        logic [WIDTH-1:0] out_1905;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1905 (
            .a(out_1902),
            .b(out_1904),
            .outp(out_1905)
        );        
        

        logic [WIDTH-1:0] out_1906;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.01626)
        ) inst_1906 (
            .outp(out_1906)
        );
        

        logic [WIDTH-1:0] out_1907;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1907 (
            .a(out_1),
            .b(out_1906),
            .outp(out_1907)
        );        
        

        logic [WIDTH-1:0] out_1908;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1908 (
            .a(out_1905),
            .b(out_1907),
            .outp(out_1908)
        );        
        

        logic [WIDTH-1:0] out_1909;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1909 (
            .a(out_1901),
            .b(out_1908),
            .outp(out_1909)
        );        
        

        logic [WIDTH-1:0] out_1910;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.27381)
        ) inst_1910 (
            .outp(out_1910)
        );
        

        logic [WIDTH-1:0] out_1911;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1911 (
            .a(out_1910),
            .b(out_1904),
            .outp(out_1911)
        );        
        

        logic [WIDTH-1:0] out_1912;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1912 (
            .a(out_1907),
            .b(out_1911),
            .outp(out_1912)
        );        
        

        logic [WIDTH-1:0] out_1913;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1913 (
            .a(out_1899),
            .b(out_1912),
            .outp(out_1913)
        );        
        

        logic [WIDTH-1:0] out_1914;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1914 (
            .a(out_1893),
            .b(out_1891),
            .outp(out_1914)
        );        
        

        logic [WIDTH-1:0] out_1915;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1915 (
            .a(out_1913),
            .b(out_1914),
            .outp(out_1915)
        );        
        

        logic [WIDTH-1:0] out_1916;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1916 (
            .a(out_1909),
            .b(out_1915),
            .outp(out_1916)
        );        
        

        logic [WIDTH-1:0] out_1917;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1917 (
            .in(out_1916),
            .outp(out_1917)
        );
        

        logic [WIDTH-1:0] out_1918;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.825)
        ) inst_1918 (
            .outp(out_1918)
        );
        

        logic [WIDTH-1:0] out_1919;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1919 (
            .a(out_1918),
            .b(out_14),
            .outp(out_1919)
        );        
        

        logic [WIDTH-1:0] out_1920;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1920 (
            .a(out_1917),
            .b(out_1919),
            .outp(out_1920)
        );        
        

        logic [WIDTH-1:0] out_1921;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.05)
        ) inst_1921 (
            .outp(out_1921)
        );
        

        logic [WIDTH-1:0] out_1922;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1922 (
            .a(out_1921),
            .b(out_14),
            .outp(out_1922)
        );        
        

        logic [WIDTH-1:0] out_1923;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1923 (
            .in(out_1922),
            .outp(out_1923)
        );
        

        logic [WIDTH-1:0] out_1924;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1924 (
            .a(out_1920),
            .b(out_1923),
            .outp(out_1924)
        );        
        

        logic [WIDTH-1:0] out_1925;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0805)
        ) inst_1925 (
            .outp(out_1925)
        );
        

        logic [WIDTH-1:0] out_1926;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1926 (
            .a(out_3),
            .b(out_1925),
            .outp(out_1926)
        );        
        

        logic [WIDTH-1:0] out_1927;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1927 (
            .a(out_1924),
            .b(out_1926),
            .outp(out_1927)
        );        
        

        logic [WIDTH-1:0] out_1928;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.9305)
        ) inst_1928 (
            .outp(out_1928)
        );
        

        logic [WIDTH-1:0] out_1929;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1929 (
            .a(out_1928),
            .b(out_3),
            .outp(out_1929)
        );        
        

        logic [WIDTH-1:0] out_1930;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1930 (
            .a(out_1927),
            .b(out_1929),
            .outp(out_1930)
        );        
        

        logic [WIDTH-1:0] out_1931;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.608333)
        ) inst_1931 (
            .outp(out_1931)
        );
        

        logic [WIDTH-1:0] out_1932;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.71003)
        ) inst_1932 (
            .outp(out_1932)
        );
        

        logic [WIDTH-1:0] out_1933;
        fixed_point_mul #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1933 (
            .a(out_13),
            .b(out_1932),
            .outp(out_1933)
        );        
        

        logic [WIDTH-1:0] out_1934;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1934 (
            .a(out_1931),
            .b(out_1933),
            .outp(out_1934)
        );        
        

        logic [WIDTH-1:0] out_1935;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1935 (
            .in(out_1934),
            .outp(out_1935)
        );
        

        logic [WIDTH-1:0] out_1936;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0055)
        ) inst_1936 (
            .outp(out_1936)
        );
        

        logic [WIDTH-1:0] out_1937;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1937 (
            .a(out_3),
            .b(out_1936),
            .outp(out_1937)
        );        
        

        logic [WIDTH-1:0] out_1938;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1938 (
            .in(out_1937),
            .outp(out_1938)
        );
        

        logic [WIDTH-1:0] out_1939;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1939 (
            .a(out_1935),
            .b(out_1938),
            .outp(out_1939)
        );        
        

        logic [WIDTH-1:0] out_1940;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1940 (
            .in(out_1939),
            .outp(out_1940)
        );
        

        logic [WIDTH-1:0] out_1941;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1941 (
            .a(out_1940),
            .b(out_460),
            .outp(out_1941)
        );        
        

        logic [WIDTH-1:0] out_1942;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1942 (
            .a(out_1930),
            .b(out_1941),
            .outp(out_1942)
        );        
        

        logic [WIDTH-1:0] out_1943;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1943 (
            .a(out_1889),
            .b(out_1942),
            .outp(out_1943)
        );        
        

        logic [WIDTH-1:0] out_1944;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1944 (
            .in(out_1919),
            .outp(out_1944)
        );
        

        logic [WIDTH-1:0] out_1945;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0305)
        ) inst_1945 (
            .outp(out_1945)
        );
        

        logic [WIDTH-1:0] out_1946;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1946 (
            .a(out_3),
            .b(out_1945),
            .outp(out_1946)
        );        
        

        logic [WIDTH-1:0] out_1947;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1947 (
            .in(out_1946),
            .outp(out_1947)
        );
        

        logic [WIDTH-1:0] out_1948;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1948 (
            .a(out_1944),
            .b(out_1947),
            .outp(out_1948)
        );        
        

        logic [WIDTH-1:0] out_1949;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1949 (
            .in(out_1948),
            .outp(out_1949)
        );
        

        logic [WIDTH-1:0] out_1950;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1950 (
            .a(out_1949),
            .b(out_460),
            .outp(out_1950)
        );        
        

        logic [WIDTH-1:0] out_1951;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1951 (
            .a(out_1943),
            .b(out_1950),
            .outp(out_1951)
        );        
        

        logic [WIDTH-1:0] out_1952;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.15)
        ) inst_1952 (
            .outp(out_1952)
        );
        

        logic [WIDTH-1:0] out_1953;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1953 (
            .a(out_1952),
            .b(out_14),
            .outp(out_1953)
        );        
        

        logic [WIDTH-1:0] out_1954;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1954 (
            .a(out_1660),
            .b(out_1953),
            .outp(out_1954)
        );        
        

        logic [WIDTH-1:0] out_1955;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.6805)
        ) inst_1955 (
            .outp(out_1955)
        );
        

        logic [WIDTH-1:0] out_1956;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1956 (
            .a(out_3),
            .b(out_1955),
            .outp(out_1956)
        );        
        

        logic [WIDTH-1:0] out_1957;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1957 (
            .a(out_1954),
            .b(out_1956),
            .outp(out_1957)
        );        
        

        logic [WIDTH-1:0] out_1958;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5805)
        ) inst_1958 (
            .outp(out_1958)
        );
        

        logic [WIDTH-1:0] out_1959;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1959 (
            .a(out_1958),
            .b(out_3),
            .outp(out_1959)
        );        
        

        logic [WIDTH-1:0] out_1960;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1960 (
            .a(out_1957),
            .b(out_1959),
            .outp(out_1960)
        );        
        

        logic [WIDTH-1:0] out_1961;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1961 (
            .a(out_1951),
            .b(out_1960),
            .outp(out_1961)
        );        
        

        logic [WIDTH-1:0] out_1962;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.8305)
        ) inst_1962 (
            .outp(out_1962)
        );
        

        logic [WIDTH-1:0] out_1963;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1963 (
            .a(out_3),
            .b(out_1962),
            .outp(out_1963)
        );        
        

        logic [WIDTH-1:0] out_1964;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1964 (
            .a(out_1675),
            .b(out_1963),
            .outp(out_1964)
        );        
        

        logic [WIDTH-1:0] out_1965;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.4305)
        ) inst_1965 (
            .outp(out_1965)
        );
        

        logic [WIDTH-1:0] out_1966;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1966 (
            .a(out_1965),
            .b(out_3),
            .outp(out_1966)
        );        
        

        logic [WIDTH-1:0] out_1967;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1967 (
            .a(out_1964),
            .b(out_1966),
            .outp(out_1967)
        );        
        

        logic [WIDTH-1:0] out_1968;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.45)
        ) inst_1968 (
            .outp(out_1968)
        );
        

        logic [WIDTH-1:0] out_1969;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1969 (
            .a(out_1968),
            .b(out_14),
            .outp(out_1969)
        );        
        

        logic [WIDTH-1:0] out_1970;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1970 (
            .in(out_1969),
            .outp(out_1970)
        );
        

        logic [WIDTH-1:0] out_1971;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1971 (
            .a(out_1967),
            .b(out_1970),
            .outp(out_1971)
        );        
        

        logic [WIDTH-1:0] out_1972;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1972 (
            .a(out_1961),
            .b(out_1971),
            .outp(out_1972)
        );        
        

        logic [WIDTH-1:0] out_1973;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1973 (
            .a(out_1860),
            .b(out_1963),
            .outp(out_1973)
        );        
        

        logic [WIDTH-1:0] out_1974;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1974 (
            .a(out_1973),
            .b(out_1966),
            .outp(out_1974)
        );        
        

        logic [WIDTH-1:0] out_1975;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1975 (
            .in(out_1953),
            .outp(out_1975)
        );
        

        logic [WIDTH-1:0] out_1976;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1976 (
            .a(out_1974),
            .b(out_1975),
            .outp(out_1976)
        );        
        

        logic [WIDTH-1:0] out_1977;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1977 (
            .in(out_1953),
            .outp(out_1977)
        );
        

        logic [WIDTH-1:0] out_1978;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1978 (
            .in(out_1963),
            .outp(out_1978)
        );
        

        logic [WIDTH-1:0] out_1979;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1979 (
            .a(out_1977),
            .b(out_1978),
            .outp(out_1979)
        );        
        

        logic [WIDTH-1:0] out_1980;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1980 (
            .in(out_1979),
            .outp(out_1980)
        );
        

        logic [WIDTH-1:0] out_1981;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1981 (
            .a(out_336),
            .b(out_1980),
            .outp(out_1981)
        );        
        

        logic [WIDTH-1:0] out_1982;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1982 (
            .a(out_1976),
            .b(out_1981),
            .outp(out_1982)
        );        
        

        logic [WIDTH-1:0] out_1983;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1983 (
            .a(out_1980),
            .b(out_343),
            .outp(out_1983)
        );        
        

        logic [WIDTH-1:0] out_1984;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1984 (
            .a(out_1982),
            .b(out_1983),
            .outp(out_1984)
        );        
        

        logic [WIDTH-1:0] out_1985;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1985 (
            .a(out_1972),
            .b(out_1984),
            .outp(out_1985)
        );        
        

        logic [WIDTH-1:0] out_1986;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.1805)
        ) inst_1986 (
            .outp(out_1986)
        );
        

        logic [WIDTH-1:0] out_1987;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1987 (
            .a(out_3),
            .b(out_1986),
            .outp(out_1987)
        );        
        

        logic [WIDTH-1:0] out_1988;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1988 (
            .a(out_1954),
            .b(out_1987),
            .outp(out_1988)
        );        
        

        logic [WIDTH-1:0] out_1989;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.0805)
        ) inst_1989 (
            .outp(out_1989)
        );
        

        logic [WIDTH-1:0] out_1990;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1990 (
            .a(out_1989),
            .b(out_3),
            .outp(out_1990)
        );        
        

        logic [WIDTH-1:0] out_1991;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1991 (
            .a(out_1988),
            .b(out_1990),
            .outp(out_1991)
        );        
        

        logic [WIDTH-1:0] out_1992;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1992 (
            .a(out_1985),
            .b(out_1991),
            .outp(out_1992)
        );        
        

        logic [WIDTH-1:0] out_1993;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1993 (
            .a(out_1752),
            .b(out_1751),
            .outp(out_1993)
        );        
        

        logic [WIDTH-1:0] out_1994;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1994 (
            .a(out_1726),
            .b(out_1993),
            .outp(out_1994)
        );        
        

        logic [WIDTH-1:0] out_1995;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1995 (
            .a(out_1748),
            .b(out_1747),
            .outp(out_1995)
        );        
        

        logic [WIDTH-1:0] out_1996;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1996 (
            .a(out_1994),
            .b(out_1995),
            .outp(out_1996)
        );        
        

        logic [WIDTH-1:0] out_1997;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1997 (
            .a(out_1992),
            .b(out_1996),
            .outp(out_1997)
        );        
        

        logic [WIDTH-1:0] out_1998;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_1998 (
            .a(out_1740),
            .b(out_1993),
            .outp(out_1998)
        );        
        

        logic [WIDTH-1:0] out_1999;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.30243)
        ) inst_1999 (
            .outp(out_1999)
        );
        

        logic [WIDTH-1:0] out_2000;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2000 (
            .a(out_1748),
            .b(out_1999),
            .outp(out_2000)
        );        
        

        logic [WIDTH-1:0] out_2001;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2001 (
            .a(out_1998),
            .b(out_2000),
            .outp(out_2001)
        );        
        

        logic [WIDTH-1:0] out_2002;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2002 (
            .a(out_1997),
            .b(out_2001),
            .outp(out_2002)
        );        
        

        logic [WIDTH-1:0] out_2003;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2003 (
            .a(out_1744),
            .b(out_1753),
            .outp(out_2003)
        );        
        

        logic [WIDTH-1:0] out_2004;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2004 (
            .a(out_1999),
            .b(out_1748),
            .outp(out_2004)
        );        
        

        logic [WIDTH-1:0] out_2005;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2005 (
            .a(out_2003),
            .b(out_2004),
            .outp(out_2005)
        );        
        

        logic [WIDTH-1:0] out_2006;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2006 (
            .a(out_2002),
            .b(out_2005),
            .outp(out_2006)
        );        
        

        logic [WIDTH-1:0] out_2007;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.2805)
        ) inst_2007 (
            .outp(out_2007)
        );
        

        logic [WIDTH-1:0] out_2008;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2008 (
            .a(out_3),
            .b(out_2007),
            .outp(out_2008)
        );        
        

        logic [WIDTH-1:0] out_2009;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2009 (
            .a(out_1676),
            .b(out_2008),
            .outp(out_2009)
        );        
        

        logic [WIDTH-1:0] out_2010;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.1805)
        ) inst_2010 (
            .outp(out_2010)
        );
        

        logic [WIDTH-1:0] out_2011;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2011 (
            .a(out_2010),
            .b(out_3),
            .outp(out_2011)
        );        
        

        logic [WIDTH-1:0] out_2012;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2012 (
            .a(out_2009),
            .b(out_2011),
            .outp(out_2012)
        );        
        

        logic [WIDTH-1:0] out_2013;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2013 (
            .a(out_2006),
            .b(out_2012),
            .outp(out_2013)
        );        
        

        logic [WIDTH-1:0] out_2014;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.52214)
        ) inst_2014 (
            .outp(out_2014)
        );
        

        logic [WIDTH-1:0] out_2015;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2015 (
            .a(out_194),
            .b(out_2014),
            .outp(out_2015)
        );        
        

        logic [WIDTH-1:0] out_2016;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2016 (
            .a(out_1676),
            .b(out_2015),
            .outp(out_2016)
        );        
        

        logic [WIDTH-1:0] out_2017;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.97215)
        ) inst_2017 (
            .outp(out_2017)
        );
        

        logic [WIDTH-1:0] out_2018;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2018 (
            .a(out_2017),
            .b(out_194),
            .outp(out_2018)
        );        
        

        logic [WIDTH-1:0] out_2019;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2019 (
            .a(out_2016),
            .b(out_2018),
            .outp(out_2019)
        );        
        

        logic [WIDTH-1:0] out_2020;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2020 (
            .in(out_1659),
            .outp(out_2020)
        );
        

        logic [WIDTH-1:0] out_2021;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.15268)
        ) inst_2021 (
            .outp(out_2021)
        );
        

        logic [WIDTH-1:0] out_2022;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2022 (
            .a(out_204),
            .b(out_2021),
            .outp(out_2022)
        );        
        

        logic [WIDTH-1:0] out_2023;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2023 (
            .in(out_2022),
            .outp(out_2023)
        );
        

        logic [WIDTH-1:0] out_2024;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2024 (
            .a(out_2020),
            .b(out_2023),
            .outp(out_2024)
        );        
        

        logic [WIDTH-1:0] out_2025;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2025 (
            .in(out_2024),
            .outp(out_2025)
        );
        

        logic [WIDTH-1:0] out_2026;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2026 (
            .a(out_200),
            .b(out_2025),
            .outp(out_2026)
        );        
        

        logic [WIDTH-1:0] out_2027;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2027 (
            .a(out_2019),
            .b(out_2026),
            .outp(out_2027)
        );        
        

        logic [WIDTH-1:0] out_2028;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2028 (
            .in(out_2015),
            .outp(out_2028)
        );
        

        logic [WIDTH-1:0] out_2029;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2029 (
            .a(out_2020),
            .b(out_2028),
            .outp(out_2029)
        );        
        

        logic [WIDTH-1:0] out_2030;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2030 (
            .in(out_2029),
            .outp(out_2030)
        );
        

        logic [WIDTH-1:0] out_2031;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2031 (
            .a(out_2030),
            .b(out_214),
            .outp(out_2031)
        );        
        

        logic [WIDTH-1:0] out_2032;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2032 (
            .a(out_2027),
            .b(out_2031),
            .outp(out_2032)
        );        
        

        logic [WIDTH-1:0] out_2033;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2033 (
            .a(out_2013),
            .b(out_2032),
            .outp(out_2033)
        );        
        

        logic [WIDTH-1:0] out_2034;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.0805)
        ) inst_2034 (
            .outp(out_2034)
        );
        

        logic [WIDTH-1:0] out_2035;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2035 (
            .a(out_3),
            .b(out_2034),
            .outp(out_2035)
        );        
        

        logic [WIDTH-1:0] out_2036;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2036 (
            .a(out_1676),
            .b(out_2035),
            .outp(out_2036)
        );        
        

        logic [WIDTH-1:0] out_2037;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.9805)
        ) inst_2037 (
            .outp(out_2037)
        );
        

        logic [WIDTH-1:0] out_2038;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2038 (
            .a(out_2037),
            .b(out_3),
            .outp(out_2038)
        );        
        

        logic [WIDTH-1:0] out_2039;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2039 (
            .a(out_2036),
            .b(out_2038),
            .outp(out_2039)
        );        
        

        logic [WIDTH-1:0] out_2040;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2040 (
            .a(out_2033),
            .b(out_2039),
            .outp(out_2040)
        );        
        

        logic [WIDTH-1:0] out_2041;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.625)
        ) inst_2041 (
            .outp(out_2041)
        );
        

        logic [WIDTH-1:0] out_2042;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2042 (
            .a(out_2041),
            .b(out_14),
            .outp(out_2042)
        );        
        

        logic [WIDTH-1:0] out_2043;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2043 (
            .in(out_2042),
            .outp(out_2043)
        );
        

        logic [WIDTH-1:0] out_2044;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2044 (
            .a(out_1675),
            .b(out_2043),
            .outp(out_2044)
        );        
        

        logic [WIDTH-1:0] out_2045;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6305)
        ) inst_2045 (
            .outp(out_2045)
        );
        

        logic [WIDTH-1:0] out_2046;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2046 (
            .a(out_3),
            .b(out_2045),
            .outp(out_2046)
        );        
        

        logic [WIDTH-1:0] out_2047;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2047 (
            .a(out_2044),
            .b(out_2046),
            .outp(out_2047)
        );        
        

        logic [WIDTH-1:0] out_2048;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.5305)
        ) inst_2048 (
            .outp(out_2048)
        );
        

        logic [WIDTH-1:0] out_2049;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2049 (
            .a(out_2048),
            .b(out_3),
            .outp(out_2049)
        );        
        

        logic [WIDTH-1:0] out_2050;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2050 (
            .a(out_2047),
            .b(out_2049),
            .outp(out_2050)
        );        
        

        logic [WIDTH-1:0] out_2051;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2051 (
            .a(out_2040),
            .b(out_2050),
            .outp(out_2051)
        );        
        

        logic [WIDTH-1:0] out_2052;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2052 (
            .a(out_1660),
            .b(out_2035),
            .outp(out_2052)
        );        
        

        logic [WIDTH-1:0] out_2053;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2053 (
            .a(out_2052),
            .b(out_2049),
            .outp(out_2053)
        );        
        

        logic [WIDTH-1:0] out_2054;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2054 (
            .a(out_2053),
            .b(out_1872),
            .outp(out_2054)
        );        
        

        logic [WIDTH-1:0] out_2055;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.8055)
        ) inst_2055 (
            .outp(out_2055)
        );
        

        logic [WIDTH-1:0] out_2056;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2056 (
            .a(out_3),
            .b(out_2055),
            .outp(out_2056)
        );        
        

        logic [WIDTH-1:0] out_2057;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2057 (
            .in(out_2056),
            .outp(out_2057)
        );
        

        logic [WIDTH-1:0] out_2058;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2058 (
            .a(out_1873),
            .b(out_2057),
            .outp(out_2058)
        );        
        

        logic [WIDTH-1:0] out_2059;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2059 (
            .in(out_2058),
            .outp(out_2059)
        );
        

        logic [WIDTH-1:0] out_2060;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2060 (
            .a(out_9),
            .b(out_2059),
            .outp(out_2060)
        );        
        

        logic [WIDTH-1:0] out_2061;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2061 (
            .a(out_2054),
            .b(out_2060),
            .outp(out_2061)
        );        
        

        logic [WIDTH-1:0] out_2062;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2062 (
            .a(out_2059),
            .b(out_21),
            .outp(out_2062)
        );        
        

        logic [WIDTH-1:0] out_2063;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2063 (
            .a(out_2061),
            .b(out_2062),
            .outp(out_2063)
        );        
        

        logic [WIDTH-1:0] out_2064;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2064 (
            .a(out_2051),
            .b(out_2063),
            .outp(out_2064)
        );        
        

        logic [WIDTH-1:0] out_2065;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0055)
        ) inst_2065 (
            .outp(out_2065)
        );
        

        logic [WIDTH-1:0] out_2066;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2066 (
            .a(out_3),
            .b(out_2065),
            .outp(out_2066)
        );        
        

        logic [WIDTH-1:0] out_2067;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2067 (
            .a(out_1870),
            .b(out_2066),
            .outp(out_2067)
        );        
        

        logic [WIDTH-1:0] out_2068;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.9055)
        ) inst_2068 (
            .outp(out_2068)
        );
        

        logic [WIDTH-1:0] out_2069;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2069 (
            .a(out_2068),
            .b(out_3),
            .outp(out_2069)
        );        
        

        logic [WIDTH-1:0] out_2070;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2070 (
            .a(out_2067),
            .b(out_2069),
            .outp(out_2070)
        );        
        

        logic [WIDTH-1:0] out_2071;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2071 (
            .a(out_2064),
            .b(out_2070),
            .outp(out_2071)
        );        
        

        logic [WIDTH-1:0] out_2072;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2072 (
            .a(out_1675),
            .b(out_1970),
            .outp(out_2072)
        );        
        

        logic [WIDTH-1:0] out_2073;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2073 (
            .a(out_2072),
            .b(out_1875),
            .outp(out_2073)
        );        
        

        logic [WIDTH-1:0] out_2074;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0055)
        ) inst_2074 (
            .outp(out_2074)
        );
        

        logic [WIDTH-1:0] out_2075;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2075 (
            .a(out_2074),
            .b(out_3),
            .outp(out_2075)
        );        
        

        logic [WIDTH-1:0] out_2076;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2076 (
            .a(out_2073),
            .b(out_2075),
            .outp(out_2076)
        );        
        

        logic [WIDTH-1:0] out_2077;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2077 (
            .a(out_2071),
            .b(out_2076),
            .outp(out_2077)
        );        
        

        logic [WIDTH-1:0] out_2078;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2078 (
            .a(out_1660),
            .b(out_1875),
            .outp(out_2078)
        );        
        

        logic [WIDTH-1:0] out_2079;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2079 (
            .a(out_2078),
            .b(out_2075),
            .outp(out_2079)
        );        
        

        logic [WIDTH-1:0] out_2080;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.8)
        ) inst_2080 (
            .outp(out_2080)
        );
        

        logic [WIDTH-1:0] out_2081;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2081 (
            .a(out_2080),
            .b(out_14),
            .outp(out_2081)
        );        
        

        logic [WIDTH-1:0] out_2082;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2082 (
            .a(out_2079),
            .b(out_2081),
            .outp(out_2082)
        );        
        

        logic [WIDTH-1:0] out_2083;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2083 (
            .a(out_2077),
            .b(out_2082),
            .outp(out_2083)
        );        
        

        logic [WIDTH-1:0] out_2084;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.57243)
        ) inst_2084 (
            .outp(out_2084)
        );
        

        logic [WIDTH-1:0] out_2085;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2085 (
            .a(out_1495),
            .b(out_2084),
            .outp(out_2085)
        );        
        

        logic [WIDTH-1:0] out_2086;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2086 (
            .a(out_3),
            .b(out_2085),
            .outp(out_2086)
        );        
        

        logic [WIDTH-1:0] out_2087;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2087 (
            .in(out_2086),
            .outp(out_2087)
        );
        

        logic [WIDTH-1:0] out_2088;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2088 (
            .a(out_753),
            .b(out_2087),
            .outp(out_2088)
        );        
        

        logic [WIDTH-1:0] out_2089;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2089 (
            .in(out_2088),
            .outp(out_2089)
        );
        

        logic [WIDTH-1:0] out_2090;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2090 (
            .a(out_9),
            .b(out_2089),
            .outp(out_2090)
        );        
        

        logic [WIDTH-1:0] out_2091;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2091 (
            .a(out_2089),
            .b(out_21),
            .outp(out_2091)
        );        
        

        logic [WIDTH-1:0] out_2092;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2092 (
            .a(out_2090),
            .b(out_2091),
            .outp(out_2092)
        );        
        

        logic [WIDTH-1:0] out_2093;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2093 (
            .a(out_2083),
            .b(out_2092),
            .outp(out_2093)
        );        
        

        logic [WIDTH-1:0] out_2094;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2094 (
            .a(out_717),
            .b(out_752),
            .outp(out_2094)
        );        
        

        logic [WIDTH-1:0] out_2095;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.051)
        ) inst_2095 (
            .outp(out_2095)
        );
        

        logic [WIDTH-1:0] out_2096;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2096 (
            .a(out_3),
            .b(out_2095),
            .outp(out_2096)
        );        
        

        logic [WIDTH-1:0] out_2097;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2097 (
            .a(out_2094),
            .b(out_2096),
            .outp(out_2097)
        );        
        

        logic [WIDTH-1:0] out_2098;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.951)
        ) inst_2098 (
            .outp(out_2098)
        );
        

        logic [WIDTH-1:0] out_2099;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2099 (
            .a(out_2098),
            .b(out_3),
            .outp(out_2099)
        );        
        

        logic [WIDTH-1:0] out_2100;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2100 (
            .a(out_2097),
            .b(out_2099),
            .outp(out_2100)
        );        
        

        logic [WIDTH-1:0] out_2101;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2101 (
            .a(out_2093),
            .b(out_2100),
            .outp(out_2101)
        );        
        

        logic [WIDTH-1:0] out_2102;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.601)
        ) inst_2102 (
            .outp(out_2102)
        );
        

        logic [WIDTH-1:0] out_2103;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2103 (
            .a(out_3),
            .b(out_2102),
            .outp(out_2103)
        );        
        

        logic [WIDTH-1:0] out_2104;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2104 (
            .a(out_718),
            .b(out_2103),
            .outp(out_2104)
        );        
        

        logic [WIDTH-1:0] out_2105;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.501)
        ) inst_2105 (
            .outp(out_2105)
        );
        

        logic [WIDTH-1:0] out_2106;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2106 (
            .a(out_2105),
            .b(out_3),
            .outp(out_2106)
        );        
        

        logic [WIDTH-1:0] out_2107;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2107 (
            .a(out_2104),
            .b(out_2106),
            .outp(out_2107)
        );        
        

        logic [WIDTH-1:0] out_2108;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2108 (
            .a(out_2101),
            .b(out_2107),
            .outp(out_2108)
        );        
        

        logic [WIDTH-1:0] out_2109;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2109 (
            .a(out_727),
            .b(out_2096),
            .outp(out_2109)
        );        
        

        logic [WIDTH-1:0] out_2110;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2110 (
            .a(out_2109),
            .b(out_2106),
            .outp(out_2110)
        );        
        

        logic [WIDTH-1:0] out_2111;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.825)
        ) inst_2111 (
            .outp(out_2111)
        );
        

        logic [WIDTH-1:0] out_2112;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2112 (
            .a(out_2111),
            .b(out_14),
            .outp(out_2112)
        );        
        

        logic [WIDTH-1:0] out_2113;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2113 (
            .in(out_2112),
            .outp(out_2113)
        );
        

        logic [WIDTH-1:0] out_2114;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2114 (
            .a(out_2110),
            .b(out_2113),
            .outp(out_2114)
        );        
        

        logic [WIDTH-1:0] out_2115;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.776)
        ) inst_2115 (
            .outp(out_2115)
        );
        

        logic [WIDTH-1:0] out_2116;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2116 (
            .a(out_3),
            .b(out_2115),
            .outp(out_2116)
        );        
        

        logic [WIDTH-1:0] out_2117;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2117 (
            .in(out_2116),
            .outp(out_2117)
        );
        

        logic [WIDTH-1:0] out_2118;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2118 (
            .a(out_753),
            .b(out_2117),
            .outp(out_2118)
        );        
        

        logic [WIDTH-1:0] out_2119;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2119 (
            .in(out_2118),
            .outp(out_2119)
        );
        

        logic [WIDTH-1:0] out_2120;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2120 (
            .a(out_9),
            .b(out_2119),
            .outp(out_2120)
        );        
        

        logic [WIDTH-1:0] out_2121;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2121 (
            .a(out_2114),
            .b(out_2120),
            .outp(out_2121)
        );        
        

        logic [WIDTH-1:0] out_2122;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2122 (
            .a(out_2119),
            .b(out_21),
            .outp(out_2122)
        );        
        

        logic [WIDTH-1:0] out_2123;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2123 (
            .a(out_2121),
            .b(out_2122),
            .outp(out_2123)
        );        
        

        logic [WIDTH-1:0] out_2124;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2124 (
            .a(out_2108),
            .b(out_2123),
            .outp(out_2124)
        );        
        

        logic [WIDTH-1:0] out_2125;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.85)
        ) inst_2125 (
            .outp(out_2125)
        );
        

        logic [WIDTH-1:0] out_2126;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2126 (
            .a(out_2125),
            .b(out_14),
            .outp(out_2126)
        );        
        

        logic [WIDTH-1:0] out_2127;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2127 (
            .in(out_2126),
            .outp(out_2127)
        );
        

        logic [WIDTH-1:0] out_2128;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2128 (
            .a(out_714),
            .b(out_2127),
            .outp(out_2128)
        );        
        

        logic [WIDTH-1:0] out_2129;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.251)
        ) inst_2129 (
            .outp(out_2129)
        );
        

        logic [WIDTH-1:0] out_2130;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2130 (
            .a(out_3),
            .b(out_2129),
            .outp(out_2130)
        );        
        

        logic [WIDTH-1:0] out_2131;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2131 (
            .a(out_2128),
            .b(out_2130),
            .outp(out_2131)
        );        
        

        logic [WIDTH-1:0] out_2132;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.151)
        ) inst_2132 (
            .outp(out_2132)
        );
        

        logic [WIDTH-1:0] out_2133;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2133 (
            .a(out_2132),
            .b(out_3),
            .outp(out_2133)
        );        
        

        logic [WIDTH-1:0] out_2134;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2134 (
            .a(out_2131),
            .b(out_2133),
            .outp(out_2134)
        );        
        

        logic [WIDTH-1:0] out_2135;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2135 (
            .a(out_2124),
            .b(out_2134),
            .outp(out_2135)
        );        
        

        logic [WIDTH-1:0] out_2136;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.45)
        ) inst_2136 (
            .outp(out_2136)
        );
        

        logic [WIDTH-1:0] out_2137;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2137 (
            .a(out_2136),
            .b(out_14),
            .outp(out_2137)
        );        
        

        logic [WIDTH-1:0] out_2138;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.55)
        ) inst_2138 (
            .outp(out_2138)
        );
        

        logic [WIDTH-1:0] out_2139;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2139 (
            .a(out_2138),
            .b(out_14),
            .outp(out_2139)
        );        
        

        logic [WIDTH-1:0] out_2140;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2140 (
            .in(out_2139),
            .outp(out_2140)
        );
        

        logic [WIDTH-1:0] out_2141;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2141 (
            .a(out_2137),
            .b(out_2140),
            .outp(out_2141)
        );        
        

        logic [WIDTH-1:0] out_2142;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.401)
        ) inst_2142 (
            .outp(out_2142)
        );
        

        logic [WIDTH-1:0] out_2143;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2143 (
            .a(out_3),
            .b(out_2142),
            .outp(out_2143)
        );        
        

        logic [WIDTH-1:0] out_2144;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2144 (
            .a(out_2141),
            .b(out_2143),
            .outp(out_2144)
        );        
        

        logic [WIDTH-1:0] out_2145;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.001)
        ) inst_2145 (
            .outp(out_2145)
        );
        

        logic [WIDTH-1:0] out_2146;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2146 (
            .a(out_2145),
            .b(out_3),
            .outp(out_2146)
        );        
        

        logic [WIDTH-1:0] out_2147;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2147 (
            .a(out_2144),
            .b(out_2146),
            .outp(out_2147)
        );        
        

        logic [WIDTH-1:0] out_2148;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2148 (
            .a(out_2135),
            .b(out_2147),
            .outp(out_2148)
        );        
        

        logic [WIDTH-1:0] out_2149;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2149 (
            .a(out_717),
            .b(out_2126),
            .outp(out_2149)
        );        
        

        logic [WIDTH-1:0] out_2150;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2150 (
            .a(out_2149),
            .b(out_2143),
            .outp(out_2150)
        );        
        

        logic [WIDTH-1:0] out_2151;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2151 (
            .a(out_2150),
            .b(out_2146),
            .outp(out_2151)
        );        
        

        logic [WIDTH-1:0] out_2152;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2152 (
            .in(out_2126),
            .outp(out_2152)
        );
        

        logic [WIDTH-1:0] out_2153;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2153 (
            .in(out_2143),
            .outp(out_2153)
        );
        

        logic [WIDTH-1:0] out_2154;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2154 (
            .a(out_2152),
            .b(out_2153),
            .outp(out_2154)
        );        
        

        logic [WIDTH-1:0] out_2155;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2155 (
            .in(out_2154),
            .outp(out_2155)
        );
        

        logic [WIDTH-1:0] out_2156;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2156 (
            .a(out_336),
            .b(out_2155),
            .outp(out_2156)
        );        
        

        logic [WIDTH-1:0] out_2157;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2157 (
            .a(out_2151),
            .b(out_2156),
            .outp(out_2157)
        );        
        

        logic [WIDTH-1:0] out_2158;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2158 (
            .a(out_2155),
            .b(out_343),
            .outp(out_2158)
        );        
        

        logic [WIDTH-1:0] out_2159;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2159 (
            .a(out_2157),
            .b(out_2158),
            .outp(out_2159)
        );        
        

        logic [WIDTH-1:0] out_2160;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2160 (
            .a(out_2148),
            .b(out_2159),
            .outp(out_2160)
        );        
        

        logic [WIDTH-1:0] out_2161;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2161 (
            .a(out_717),
            .b(out_727),
            .outp(out_2161)
        );        
        

        logic [WIDTH-1:0] out_2162;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.943)
        ) inst_2162 (
            .outp(out_2162)
        );
        

        logic [WIDTH-1:0] out_2163;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2163 (
            .a(out_3),
            .b(out_2162),
            .outp(out_2163)
        );        
        

        logic [WIDTH-1:0] out_2164;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2164 (
            .a(out_2161),
            .b(out_2163),
            .outp(out_2164)
        );        
        

        logic [WIDTH-1:0] out_2165;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.843)
        ) inst_2165 (
            .outp(out_2165)
        );
        

        logic [WIDTH-1:0] out_2166;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2166 (
            .a(out_2165),
            .b(out_3),
            .outp(out_2166)
        );        
        

        logic [WIDTH-1:0] out_2167;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2167 (
            .a(out_2164),
            .b(out_2166),
            .outp(out_2167)
        );        
        

        logic [WIDTH-1:0] out_2168;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2168 (
            .a(out_2160),
            .b(out_2167),
            .outp(out_2168)
        );        
        

        logic [WIDTH-1:0] out_2169;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.18286)
        ) inst_2169 (
            .outp(out_2169)
        );
        

        logic [WIDTH-1:0] out_2170;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2170 (
            .a(out_194),
            .b(out_2169),
            .outp(out_2170)
        );        
        

        logic [WIDTH-1:0] out_2171;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2171 (
            .a(out_2161),
            .b(out_2170),
            .outp(out_2171)
        );        
        

        logic [WIDTH-1:0] out_2172;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.63286)
        ) inst_2172 (
            .outp(out_2172)
        );
        

        logic [WIDTH-1:0] out_2173;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2173 (
            .a(out_2172),
            .b(out_194),
            .outp(out_2173)
        );        
        

        logic [WIDTH-1:0] out_2174;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2174 (
            .a(out_2171),
            .b(out_2173),
            .outp(out_2174)
        );        
        

        logic [WIDTH-1:0] out_2175;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2175 (
            .in(out_716),
            .outp(out_2175)
        );
        

        logic [WIDTH-1:0] out_2176;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.97857)
        ) inst_2176 (
            .outp(out_2176)
        );
        

        logic [WIDTH-1:0] out_2177;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2177 (
            .a(out_204),
            .b(out_2176),
            .outp(out_2177)
        );        
        

        logic [WIDTH-1:0] out_2178;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2178 (
            .in(out_2177),
            .outp(out_2178)
        );
        

        logic [WIDTH-1:0] out_2179;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2179 (
            .a(out_2175),
            .b(out_2178),
            .outp(out_2179)
        );        
        

        logic [WIDTH-1:0] out_2180;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2180 (
            .in(out_2179),
            .outp(out_2180)
        );
        

        logic [WIDTH-1:0] out_2181;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2181 (
            .a(out_200),
            .b(out_2180),
            .outp(out_2181)
        );        
        

        logic [WIDTH-1:0] out_2182;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2182 (
            .a(out_2174),
            .b(out_2181),
            .outp(out_2182)
        );        
        

        logic [WIDTH-1:0] out_2183;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2183 (
            .in(out_2170),
            .outp(out_2183)
        );
        

        logic [WIDTH-1:0] out_2184;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2184 (
            .a(out_2175),
            .b(out_2183),
            .outp(out_2184)
        );        
        

        logic [WIDTH-1:0] out_2185;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2185 (
            .in(out_2184),
            .outp(out_2185)
        );
        

        logic [WIDTH-1:0] out_2186;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2186 (
            .a(out_2185),
            .b(out_214),
            .outp(out_2186)
        );        
        

        logic [WIDTH-1:0] out_2187;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2187 (
            .a(out_2182),
            .b(out_2186),
            .outp(out_2187)
        );        
        

        logic [WIDTH-1:0] out_2188;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2188 (
            .a(out_2168),
            .b(out_2187),
            .outp(out_2188)
        );        
        

        logic [WIDTH-1:0] out_2189;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.981)
        ) inst_2189 (
            .outp(out_2189)
        );
        

        logic [WIDTH-1:0] out_2190;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2190 (
            .a(out_3),
            .b(out_2189),
            .outp(out_2190)
        );        
        

        logic [WIDTH-1:0] out_2191;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2191 (
            .a(out_2161),
            .b(out_2190),
            .outp(out_2191)
        );        
        

        logic [WIDTH-1:0] out_2192;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.881)
        ) inst_2192 (
            .outp(out_2192)
        );
        

        logic [WIDTH-1:0] out_2193;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2193 (
            .a(out_2192),
            .b(out_3),
            .outp(out_2193)
        );        
        

        logic [WIDTH-1:0] out_2194;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2194 (
            .a(out_2191),
            .b(out_2193),
            .outp(out_2194)
        );        
        

        logic [WIDTH-1:0] out_2195;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2195 (
            .a(out_2188),
            .b(out_2194),
            .outp(out_2195)
        );        
        

        logic [WIDTH-1:0] out_2196;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.4)
        ) inst_2196 (
            .outp(out_2196)
        );
        

        logic [WIDTH-1:0] out_2197;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2197 (
            .a(out_2196),
            .b(out_14),
            .outp(out_2197)
        );        
        

        logic [WIDTH-1:0] out_2198;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2198 (
            .in(out_2197),
            .outp(out_2198)
        );
        

        logic [WIDTH-1:0] out_2199;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.931)
        ) inst_2199 (
            .outp(out_2199)
        );
        

        logic [WIDTH-1:0] out_2200;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2200 (
            .a(out_3),
            .b(out_2199),
            .outp(out_2200)
        );        
        

        logic [WIDTH-1:0] out_2201;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2201 (
            .in(out_2200),
            .outp(out_2201)
        );
        

        logic [WIDTH-1:0] out_2202;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2202 (
            .a(out_2198),
            .b(out_2201),
            .outp(out_2202)
        );        
        

        logic [WIDTH-1:0] out_2203;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2203 (
            .in(out_2202),
            .outp(out_2203)
        );
        

        logic [WIDTH-1:0] out_2204;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2204 (
            .a(out_2203),
            .b(out_460),
            .outp(out_2204)
        );        
        

        logic [WIDTH-1:0] out_2205;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2205 (
            .a(out_2195),
            .b(out_2204),
            .outp(out_2205)
        );        
        

        logic [WIDTH-1:0] out_2206;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.656)
        ) inst_2206 (
            .outp(out_2206)
        );
        

        logic [WIDTH-1:0] out_2207;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2207 (
            .a(out_2206),
            .b(out_3),
            .outp(out_2207)
        );        
        

        logic [WIDTH-1:0] out_2208;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2208 (
            .a(out_718),
            .b(out_2207),
            .outp(out_2208)
        );        
        

        logic [WIDTH-1:0] out_2209;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.756)
        ) inst_2209 (
            .outp(out_2209)
        );
        

        logic [WIDTH-1:0] out_2210;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2210 (
            .a(out_3),
            .b(out_2209),
            .outp(out_2210)
        );        
        

        logic [WIDTH-1:0] out_2211;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2211 (
            .a(out_2208),
            .b(out_2210),
            .outp(out_2211)
        );        
        

        logic [WIDTH-1:0] out_2212;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2212 (
            .a(out_2205),
            .b(out_2211),
            .outp(out_2212)
        );        
        

        logic [WIDTH-1:0] out_2213;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.48101)
        ) inst_2213 (
            .outp(out_2213)
        );
        

        logic [WIDTH-1:0] out_2214;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2214 (
            .a(out_2213),
            .b(out_3),
            .outp(out_2214)
        );        
        

        logic [WIDTH-1:0] out_2215;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2215 (
            .a(out_731),
            .b(out_2214),
            .outp(out_2215)
        );        
        

        logic [WIDTH-1:0] out_2216;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.656)
        ) inst_2216 (
            .outp(out_2216)
        );
        

        logic [WIDTH-1:0] out_2217;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2217 (
            .a(out_3),
            .b(out_2216),
            .outp(out_2217)
        );        
        

        logic [WIDTH-1:0] out_2218;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2218 (
            .a(out_2215),
            .b(out_2217),
            .outp(out_2218)
        );        
        

        logic [WIDTH-1:0] out_2219;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2219 (
            .a(out_2212),
            .b(out_2218),
            .outp(out_2219)
        );        
        

        logic [WIDTH-1:0] out_2220;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2220 (
            .a(out_717),
            .b(out_742),
            .outp(out_2220)
        );        
        

        logic [WIDTH-1:0] out_2221;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2221 (
            .a(out_2220),
            .b(out_2214),
            .outp(out_2221)
        );        
        

        logic [WIDTH-1:0] out_2222;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2222 (
            .a(out_2221),
            .b(out_2217),
            .outp(out_2222)
        );        
        

        logic [WIDTH-1:0] out_2223;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2223 (
            .a(out_2219),
            .b(out_2222),
            .outp(out_2223)
        );        
        

        logic [WIDTH-1:0] out_2224;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.756)
        ) inst_2224 (
            .outp(out_2224)
        );
        

        logic [WIDTH-1:0] out_2225;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2225 (
            .a(out_2224),
            .b(out_3),
            .outp(out_2225)
        );        
        

        logic [WIDTH-1:0] out_2226;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2226 (
            .a(out_718),
            .b(out_2225),
            .outp(out_2226)
        );        
        

        logic [WIDTH-1:0] out_2227;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.481)
        ) inst_2227 (
            .outp(out_2227)
        );
        

        logic [WIDTH-1:0] out_2228;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2228 (
            .a(out_3),
            .b(out_2227),
            .outp(out_2228)
        );        
        

        logic [WIDTH-1:0] out_2229;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2229 (
            .a(out_2226),
            .b(out_2228),
            .outp(out_2229)
        );        
        

        logic [WIDTH-1:0] out_2230;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2230 (
            .in(out_2214),
            .outp(out_2230)
        );
        

        logic [WIDTH-1:0] out_2231;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2231 (
            .a(out_753),
            .b(out_2230),
            .outp(out_2231)
        );        
        

        logic [WIDTH-1:0] out_2232;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2232 (
            .in(out_2231),
            .outp(out_2232)
        );
        

        logic [WIDTH-1:0] out_2233;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2233 (
            .a(out_9),
            .b(out_2232),
            .outp(out_2233)
        );        
        

        logic [WIDTH-1:0] out_2234;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2234 (
            .a(out_2229),
            .b(out_2233),
            .outp(out_2234)
        );        
        

        logic [WIDTH-1:0] out_2235;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2235 (
            .a(out_2232),
            .b(out_21),
            .outp(out_2235)
        );        
        

        logic [WIDTH-1:0] out_2236;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2236 (
            .a(out_2234),
            .b(out_2235),
            .outp(out_2236)
        );        
        

        logic [WIDTH-1:0] out_2237;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2237 (
            .a(out_2223),
            .b(out_2236),
            .outp(out_2237)
        );        
        

        logic [WIDTH-1:0] out_2238;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.775)
        ) inst_2238 (
            .outp(out_2238)
        );
        

        logic [WIDTH-1:0] out_2239;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2239 (
            .a(out_2238),
            .b(out_14),
            .outp(out_2239)
        );        
        

        logic [WIDTH-1:0] out_2240;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2240 (
            .a(out_717),
            .b(out_2239),
            .outp(out_2240)
        );        
        

        logic [WIDTH-1:0] out_2241;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.431)
        ) inst_2241 (
            .outp(out_2241)
        );
        

        logic [WIDTH-1:0] out_2242;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2242 (
            .a(out_3),
            .b(out_2241),
            .outp(out_2242)
        );        
        

        logic [WIDTH-1:0] out_2243;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2243 (
            .a(out_2240),
            .b(out_2242),
            .outp(out_2243)
        );        
        

        logic [WIDTH-1:0] out_2244;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.331)
        ) inst_2244 (
            .outp(out_2244)
        );
        

        logic [WIDTH-1:0] out_2245;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2245 (
            .a(out_2244),
            .b(out_3),
            .outp(out_2245)
        );        
        

        logic [WIDTH-1:0] out_2246;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2246 (
            .a(out_2243),
            .b(out_2245),
            .outp(out_2246)
        );        
        

        logic [WIDTH-1:0] out_2247;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2247 (
            .a(out_2237),
            .b(out_2246),
            .outp(out_2247)
        );        
        

        logic [WIDTH-1:0] out_2248;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.981)
        ) inst_2248 (
            .outp(out_2248)
        );
        

        logic [WIDTH-1:0] out_2249;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2249 (
            .a(out_3),
            .b(out_2248),
            .outp(out_2249)
        );        
        

        logic [WIDTH-1:0] out_2250;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2250 (
            .a(out_2161),
            .b(out_2249),
            .outp(out_2250)
        );        
        

        logic [WIDTH-1:0] out_2251;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.881)
        ) inst_2251 (
            .outp(out_2251)
        );
        

        logic [WIDTH-1:0] out_2252;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2252 (
            .a(out_2251),
            .b(out_3),
            .outp(out_2252)
        );        
        

        logic [WIDTH-1:0] out_2253;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2253 (
            .a(out_2250),
            .b(out_2252),
            .outp(out_2253)
        );        
        

        logic [WIDTH-1:0] out_2254;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2254 (
            .a(out_2247),
            .b(out_2253),
            .outp(out_2254)
        );        
        

        logic [WIDTH-1:0] out_2255;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2255 (
            .a(out_727),
            .b(out_2242),
            .outp(out_2255)
        );        
        

        logic [WIDTH-1:0] out_2256;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2256 (
            .a(out_2255),
            .b(out_2252),
            .outp(out_2256)
        );        
        

        logic [WIDTH-1:0] out_2257;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.775)
        ) inst_2257 (
            .outp(out_2257)
        );
        

        logic [WIDTH-1:0] out_2258;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2258 (
            .a(out_2257),
            .b(out_14),
            .outp(out_2258)
        );        
        

        logic [WIDTH-1:0] out_2259;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2259 (
            .in(out_2258),
            .outp(out_2259)
        );
        

        logic [WIDTH-1:0] out_2260;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2260 (
            .a(out_2256),
            .b(out_2259),
            .outp(out_2260)
        );        
        

        logic [WIDTH-1:0] out_2261;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.156)
        ) inst_2261 (
            .outp(out_2261)
        );
        

        logic [WIDTH-1:0] out_2262;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2262 (
            .a(out_3),
            .b(out_2261),
            .outp(out_2262)
        );        
        

        logic [WIDTH-1:0] out_2263;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2263 (
            .in(out_2262),
            .outp(out_2263)
        );
        

        logic [WIDTH-1:0] out_2264;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2264 (
            .a(out_753),
            .b(out_2263),
            .outp(out_2264)
        );        
        

        logic [WIDTH-1:0] out_2265;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2265 (
            .in(out_2264),
            .outp(out_2265)
        );
        

        logic [WIDTH-1:0] out_2266;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2266 (
            .a(out_9),
            .b(out_2265),
            .outp(out_2266)
        );        
        

        logic [WIDTH-1:0] out_2267;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2267 (
            .a(out_2260),
            .b(out_2266),
            .outp(out_2267)
        );        
        

        logic [WIDTH-1:0] out_2268;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2268 (
            .a(out_2265),
            .b(out_21),
            .outp(out_2268)
        );        
        

        logic [WIDTH-1:0] out_2269;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2269 (
            .a(out_2267),
            .b(out_2268),
            .outp(out_2269)
        );        
        

        logic [WIDTH-1:0] out_2270;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2270 (
            .a(out_2254),
            .b(out_2269),
            .outp(out_2270)
        );        
        

        logic [WIDTH-1:0] out_2271;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.75)
        ) inst_2271 (
            .outp(out_2271)
        );
        

        logic [WIDTH-1:0] out_2272;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2272 (
            .a(out_2271),
            .b(out_14),
            .outp(out_2272)
        );        
        

        logic [WIDTH-1:0] out_2273;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2273 (
            .a(out_717),
            .b(out_2272),
            .outp(out_2273)
        );        
        

        logic [WIDTH-1:0] out_2274;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.761)
        ) inst_2274 (
            .outp(out_2274)
        );
        

        logic [WIDTH-1:0] out_2275;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2275 (
            .a(out_3),
            .b(out_2274),
            .outp(out_2275)
        );        
        

        logic [WIDTH-1:0] out_2276;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2276 (
            .a(out_2273),
            .b(out_2275),
            .outp(out_2276)
        );        
        

        logic [WIDTH-1:0] out_2277;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.661)
        ) inst_2277 (
            .outp(out_2277)
        );
        

        logic [WIDTH-1:0] out_2278;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2278 (
            .a(out_2277),
            .b(out_3),
            .outp(out_2278)
        );        
        

        logic [WIDTH-1:0] out_2279;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2279 (
            .a(out_2276),
            .b(out_2278),
            .outp(out_2279)
        );        
        

        logic [WIDTH-1:0] out_2280;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2280 (
            .a(out_2270),
            .b(out_2279),
            .outp(out_2280)
        );        
        

        logic [WIDTH-1:0] out_2281;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.167999)
        ) inst_2281 (
            .outp(out_2281)
        );
        

        logic [WIDTH-1:0] out_2282;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2282 (
            .a(out_3),
            .b(out_2281),
            .outp(out_2282)
        );        
        

        logic [WIDTH-1:0] out_2283;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2283 (
            .in(out_2282),
            .outp(out_2283)
        );
        

        logic [WIDTH-1:0] out_2284;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2284 (
            .a(out_753),
            .b(out_2283),
            .outp(out_2284)
        );        
        

        logic [WIDTH-1:0] out_2285;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2285 (
            .in(out_2284),
            .outp(out_2285)
        );
        

        logic [WIDTH-1:0] out_2286;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2286 (
            .a(out_9),
            .b(out_2285),
            .outp(out_2286)
        );        
        

        logic [WIDTH-1:0] out_2287;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2287 (
            .a(out_2285),
            .b(out_21),
            .outp(out_2287)
        );        
        

        logic [WIDTH-1:0] out_2288;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2288 (
            .a(out_2286),
            .b(out_2287),
            .outp(out_2288)
        );        
        

        logic [WIDTH-1:0] out_2289;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.48625)
        ) inst_2289 (
            .outp(out_2289)
        );
        

        logic [WIDTH-1:0] out_2290;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2290 (
            .a(out_2289),
            .b(out_553),
            .outp(out_2290)
        );        
        

        logic [WIDTH-1:0] out_2291;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.750575)
        ) inst_2291 (
            .outp(out_2291)
        );
        

        logic [WIDTH-1:0] out_2292;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2292 (
            .a(out_2291),
            .b(out_559),
            .outp(out_2292)
        );        
        

        logic [WIDTH-1:0] out_2293;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2293 (
            .a(out_556),
            .b(out_2292),
            .outp(out_2293)
        );        
        

        logic [WIDTH-1:0] out_2294;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2294 (
            .a(out_2290),
            .b(out_2293),
            .outp(out_2294)
        );        
        

        logic [WIDTH-1:0] out_2295;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.91443)
        ) inst_2295 (
            .outp(out_2295)
        );
        

        logic [WIDTH-1:0] out_2296;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2296 (
            .a(out_2295),
            .b(out_556),
            .outp(out_2296)
        );        
        

        logic [WIDTH-1:0] out_2297;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2297 (
            .a(out_2296),
            .b(out_566),
            .outp(out_2297)
        );        
        

        logic [WIDTH-1:0] out_2298;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2298 (
            .in(out_2297),
            .outp(out_2298)
        );
        

        logic [WIDTH-1:0] out_2299;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2299 (
            .a(out_2294),
            .b(out_2298),
            .outp(out_2299)
        );        
        

        logic [WIDTH-1:0] out_2300;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2300 (
            .in(out_2290),
            .outp(out_2300)
        );
        

        logic [WIDTH-1:0] out_2301;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.91443)
        ) inst_2301 (
            .outp(out_2301)
        );
        

        logic [WIDTH-1:0] out_2302;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2302 (
            .a(out_2301),
            .b(out_556),
            .outp(out_2302)
        );        
        

        logic [WIDTH-1:0] out_2303;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2303 (
            .a(out_2302),
            .b(out_566),
            .outp(out_2303)
        );        
        

        logic [WIDTH-1:0] out_2304;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2304 (
            .a(out_2300),
            .b(out_2303),
            .outp(out_2304)
        );        
        

        logic [WIDTH-1:0] out_2305;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2305 (
            .a(out_2292),
            .b(out_556),
            .outp(out_2305)
        );        
        

        logic [WIDTH-1:0] out_2306;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2306 (
            .a(out_2304),
            .b(out_2305),
            .outp(out_2306)
        );        
        

        logic [WIDTH-1:0] out_2307;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2307 (
            .a(out_2299),
            .b(out_2306),
            .outp(out_2307)
        );        
        

        logic [WIDTH-1:0] out_2308;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2308 (
            .in(out_2307),
            .outp(out_2308)
        );
        

        logic [WIDTH-1:0] out_2309;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2309 (
            .a(out_2288),
            .b(out_2308),
            .outp(out_2309)
        );        
        

        logic [WIDTH-1:0] out_2310;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.785)
        ) inst_2310 (
            .outp(out_2310)
        );
        

        logic [WIDTH-1:0] out_2311;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2311 (
            .a(out_2310),
            .b(out_14),
            .outp(out_2311)
        );        
        

        logic [WIDTH-1:0] out_2312;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.875)
        ) inst_2312 (
            .outp(out_2312)
        );
        

        logic [WIDTH-1:0] out_2313;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2313 (
            .a(out_2312),
            .b(out_14),
            .outp(out_2313)
        );        
        

        logic [WIDTH-1:0] out_2314;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2314 (
            .in(out_2313),
            .outp(out_2314)
        );
        

        logic [WIDTH-1:0] out_2315;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2315 (
            .a(out_2311),
            .b(out_2314),
            .outp(out_2315)
        );        
        

        logic [WIDTH-1:0] out_2316;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.443)
        ) inst_2316 (
            .outp(out_2316)
        );
        

        logic [WIDTH-1:0] out_2317;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2317 (
            .a(out_3),
            .b(out_2316),
            .outp(out_2317)
        );        
        

        logic [WIDTH-1:0] out_2318;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2318 (
            .a(out_2315),
            .b(out_2317),
            .outp(out_2318)
        );        
        

        logic [WIDTH-1:0] out_2319;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0570004)
        ) inst_2319 (
            .outp(out_2319)
        );
        

        logic [WIDTH-1:0] out_2320;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2320 (
            .a(out_2319),
            .b(out_3),
            .outp(out_2320)
        );        
        

        logic [WIDTH-1:0] out_2321;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2321 (
            .in(out_2320),
            .outp(out_2321)
        );
        

        logic [WIDTH-1:0] out_2322;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2322 (
            .a(out_2318),
            .b(out_2321),
            .outp(out_2322)
        );        
        

        logic [WIDTH-1:0] out_2323;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2323 (
            .a(out_2309),
            .b(out_2322),
            .outp(out_2323)
        );        
        

        logic [WIDTH-1:0] out_2324;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2324 (
            .a(out_2323),
            .b(out_2287),
            .outp(out_2324)
        );        
        

        logic [WIDTH-1:0] out_2325;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2325 (
            .a(out_2280),
            .b(out_2324),
            .outp(out_2325)
        );        
        

        logic [WIDTH-1:0] out_2326;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.207)
        ) inst_2326 (
            .outp(out_2326)
        );
        

        logic [WIDTH-1:0] out_2327;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2327 (
            .a(out_2326),
            .b(out_3),
            .outp(out_2327)
        );        
        

        logic [WIDTH-1:0] out_2328;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.707)
        ) inst_2328 (
            .outp(out_2328)
        );
        

        logic [WIDTH-1:0] out_2329;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2329 (
            .a(out_2328),
            .b(out_3),
            .outp(out_2329)
        );        
        

        logic [WIDTH-1:0] out_2330;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2330 (
            .in(out_2329),
            .outp(out_2330)
        );
        

        logic [WIDTH-1:0] out_2331;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2331 (
            .a(out_2327),
            .b(out_2330),
            .outp(out_2331)
        );        
        

        logic [WIDTH-1:0] out_2332;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2332 (
            .a(out_2331),
            .b(out_2311),
            .outp(out_2332)
        );        
        

        logic [WIDTH-1:0] out_2333;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2333 (
            .a(out_2332),
            .b(out_2314),
            .outp(out_2333)
        );        
        

        logic [WIDTH-1:0] out_2334;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.482)
        ) inst_2334 (
            .outp(out_2334)
        );
        

        logic [WIDTH-1:0] out_2335;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2335 (
            .a(out_2334),
            .b(out_3),
            .outp(out_2335)
        );        
        

        logic [WIDTH-1:0] out_2336;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2336 (
            .in(out_2335),
            .outp(out_2336)
        );
        

        logic [WIDTH-1:0] out_2337;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2337 (
            .a(out_753),
            .b(out_2336),
            .outp(out_2337)
        );        
        

        logic [WIDTH-1:0] out_2338;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2338 (
            .in(out_2337),
            .outp(out_2338)
        );
        

        logic [WIDTH-1:0] out_2339;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2339 (
            .a(out_2338),
            .b(out_21),
            .outp(out_2339)
        );        
        

        logic [WIDTH-1:0] out_2340;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.571825)
        ) inst_2340 (
            .outp(out_2340)
        );
        

        logic [WIDTH-1:0] out_2341;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2341 (
            .a(out_2340),
            .b(out_559),
            .outp(out_2341)
        );        
        

        logic [WIDTH-1:0] out_2342;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2342 (
            .a(out_556),
            .b(out_2341),
            .outp(out_2342)
        );        
        

        logic [WIDTH-1:0] out_2343;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.09318)
        ) inst_2343 (
            .outp(out_2343)
        );
        

        logic [WIDTH-1:0] out_2344;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2344 (
            .a(out_2343),
            .b(out_556),
            .outp(out_2344)
        );        
        

        logic [WIDTH-1:0] out_2345;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2345 (
            .a(out_2344),
            .b(out_566),
            .outp(out_2345)
        );        
        

        logic [WIDTH-1:0] out_2346;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2346 (
            .in(out_2345),
            .outp(out_2346)
        );
        

        logic [WIDTH-1:0] out_2347;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2347 (
            .a(out_2342),
            .b(out_2346),
            .outp(out_2347)
        );        
        

        logic [WIDTH-1:0] out_2348;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2348 (
            .a(out_2347),
            .b(out_2290),
            .outp(out_2348)
        );        
        

        logic [WIDTH-1:0] out_2349;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2349 (
            .a(out_2341),
            .b(out_556),
            .outp(out_2349)
        );        
        

        logic [WIDTH-1:0] out_2350;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2350 (
            .a(out_2345),
            .b(out_2349),
            .outp(out_2350)
        );        
        

        logic [WIDTH-1:0] out_2351;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2351 (
            .a(out_2350),
            .b(out_2300),
            .outp(out_2351)
        );        
        

        logic [WIDTH-1:0] out_2352;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2352 (
            .a(out_2348),
            .b(out_2351),
            .outp(out_2352)
        );        
        

        logic [WIDTH-1:0] out_2353;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2353 (
            .in(out_2352),
            .outp(out_2353)
        );
        

        logic [WIDTH-1:0] out_2354;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2354 (
            .a(out_2339),
            .b(out_2353),
            .outp(out_2354)
        );        
        

        logic [WIDTH-1:0] out_2355;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2355 (
            .a(out_9),
            .b(out_2338),
            .outp(out_2355)
        );        
        

        logic [WIDTH-1:0] out_2356;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2356 (
            .a(out_2354),
            .b(out_2355),
            .outp(out_2356)
        );        
        

        logic [WIDTH-1:0] out_2357;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2357 (
            .a(out_2333),
            .b(out_2356),
            .outp(out_2357)
        );        
        

        logic [WIDTH-1:0] out_2358;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2358 (
            .a(out_2339),
            .b(out_2357),
            .outp(out_2358)
        );        
        

        logic [WIDTH-1:0] out_2359;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2359 (
            .a(out_2325),
            .b(out_2358),
            .outp(out_2359)
        );        
        

        logic [WIDTH-1:0] out_2360;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.957)
        ) inst_2360 (
            .outp(out_2360)
        );
        

        logic [WIDTH-1:0] out_2361;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2361 (
            .a(out_2360),
            .b(out_3),
            .outp(out_2361)
        );        
        

        logic [WIDTH-1:0] out_2362;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2362 (
            .in(out_2361),
            .outp(out_2362)
        );
        

        logic [WIDTH-1:0] out_2363;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2363 (
            .a(out_718),
            .b(out_2362),
            .outp(out_2363)
        );        
        

        logic [WIDTH-1:0] out_2364;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.857)
        ) inst_2364 (
            .outp(out_2364)
        );
        

        logic [WIDTH-1:0] out_2365;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2365 (
            .a(out_2364),
            .b(out_3),
            .outp(out_2365)
        );        
        

        logic [WIDTH-1:0] out_2366;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2366 (
            .a(out_2363),
            .b(out_2365),
            .outp(out_2366)
        );        
        

        logic [WIDTH-1:0] out_2367;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2367 (
            .a(out_2359),
            .b(out_2366),
            .outp(out_2367)
        );        
        

        logic [WIDTH-1:0] out_2368;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.132)
        ) inst_2368 (
            .outp(out_2368)
        );
        

        logic [WIDTH-1:0] out_2369;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2369 (
            .a(out_2368),
            .b(out_3),
            .outp(out_2369)
        );        
        

        logic [WIDTH-1:0] out_2370;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2370 (
            .in(out_2369),
            .outp(out_2370)
        );
        

        logic [WIDTH-1:0] out_2371;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2371 (
            .a(out_731),
            .b(out_2370),
            .outp(out_2371)
        );        
        

        logic [WIDTH-1:0] out_2372;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.957)
        ) inst_2372 (
            .outp(out_2372)
        );
        

        logic [WIDTH-1:0] out_2373;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2373 (
            .a(out_2372),
            .b(out_3),
            .outp(out_2373)
        );        
        

        logic [WIDTH-1:0] out_2374;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2374 (
            .a(out_2371),
            .b(out_2373),
            .outp(out_2374)
        );        
        

        logic [WIDTH-1:0] out_2375;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2375 (
            .a(out_2367),
            .b(out_2374),
            .outp(out_2375)
        );        
        

        logic [WIDTH-1:0] out_2376;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2376 (
            .a(out_2220),
            .b(out_2370),
            .outp(out_2376)
        );        
        

        logic [WIDTH-1:0] out_2377;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2377 (
            .a(out_2376),
            .b(out_2373),
            .outp(out_2377)
        );        
        

        logic [WIDTH-1:0] out_2378;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2378 (
            .a(out_2375),
            .b(out_2377),
            .outp(out_2378)
        );        
        

        logic [WIDTH-1:0] out_2379;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.857)
        ) inst_2379 (
            .outp(out_2379)
        );
        

        logic [WIDTH-1:0] out_2380;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2380 (
            .a(out_2379),
            .b(out_3),
            .outp(out_2380)
        );        
        

        logic [WIDTH-1:0] out_2381;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2381 (
            .in(out_2380),
            .outp(out_2381)
        );
        

        logic [WIDTH-1:0] out_2382;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2382 (
            .a(out_718),
            .b(out_2381),
            .outp(out_2382)
        );        
        

        logic [WIDTH-1:0] out_2383;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.132)
        ) inst_2383 (
            .outp(out_2383)
        );
        

        logic [WIDTH-1:0] out_2384;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2384 (
            .a(out_2383),
            .b(out_3),
            .outp(out_2384)
        );        
        

        logic [WIDTH-1:0] out_2385;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2385 (
            .a(out_2382),
            .b(out_2384),
            .outp(out_2385)
        );        
        

        logic [WIDTH-1:0] out_2386;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2386 (
            .in(out_2370),
            .outp(out_2386)
        );
        

        logic [WIDTH-1:0] out_2387;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2387 (
            .a(out_753),
            .b(out_2386),
            .outp(out_2387)
        );        
        

        logic [WIDTH-1:0] out_2388;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2388 (
            .in(out_2387),
            .outp(out_2388)
        );
        

        logic [WIDTH-1:0] out_2389;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2389 (
            .a(out_9),
            .b(out_2388),
            .outp(out_2389)
        );        
        

        logic [WIDTH-1:0] out_2390;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2390 (
            .a(out_2385),
            .b(out_2389),
            .outp(out_2390)
        );        
        

        logic [WIDTH-1:0] out_2391;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2391 (
            .a(out_2388),
            .b(out_21),
            .outp(out_2391)
        );        
        

        logic [WIDTH-1:0] out_2392;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2392 (
            .a(out_2390),
            .b(out_2391),
            .outp(out_2392)
        );        
        

        logic [WIDTH-1:0] out_2393;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2393 (
            .a(out_2378),
            .b(out_2392),
            .outp(out_2393)
        );        
        

        logic [WIDTH-1:0] out_2394;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.282)
        ) inst_2394 (
            .outp(out_2394)
        );
        

        logic [WIDTH-1:0] out_2395;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2395 (
            .a(out_2394),
            .b(out_3),
            .outp(out_2395)
        );        
        

        logic [WIDTH-1:0] out_2396;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2396 (
            .in(out_2395),
            .outp(out_2396)
        );
        

        logic [WIDTH-1:0] out_2397;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2397 (
            .a(out_718),
            .b(out_2396),
            .outp(out_2397)
        );        
        

        logic [WIDTH-1:0] out_2398;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.182)
        ) inst_2398 (
            .outp(out_2398)
        );
        

        logic [WIDTH-1:0] out_2399;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2399 (
            .a(out_2398),
            .b(out_3),
            .outp(out_2399)
        );        
        

        logic [WIDTH-1:0] out_2400;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2400 (
            .a(out_2397),
            .b(out_2399),
            .outp(out_2400)
        );        
        

        logic [WIDTH-1:0] out_2401;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2401 (
            .a(out_2393),
            .b(out_2400),
            .outp(out_2401)
        );        
        

        logic [WIDTH-1:0] out_2402;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2402 (
            .a(out_731),
            .b(out_2395),
            .outp(out_2402)
        );        
        

        logic [WIDTH-1:0] out_2403;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.457)
        ) inst_2403 (
            .outp(out_2403)
        );
        

        logic [WIDTH-1:0] out_2404;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2404 (
            .a(out_2403),
            .b(out_3),
            .outp(out_2404)
        );        
        

        logic [WIDTH-1:0] out_2405;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2405 (
            .in(out_2404),
            .outp(out_2405)
        );
        

        logic [WIDTH-1:0] out_2406;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2406 (
            .a(out_2402),
            .b(out_2405),
            .outp(out_2406)
        );        
        

        logic [WIDTH-1:0] out_2407;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2407 (
            .a(out_2401),
            .b(out_2406),
            .outp(out_2407)
        );        
        

        logic [WIDTH-1:0] out_2408;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2408 (
            .a(out_2220),
            .b(out_2395),
            .outp(out_2408)
        );        
        

        logic [WIDTH-1:0] out_2409;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2409 (
            .a(out_2408),
            .b(out_2405),
            .outp(out_2409)
        );        
        

        logic [WIDTH-1:0] out_2410;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2410 (
            .a(out_2407),
            .b(out_2409),
            .outp(out_2410)
        );        
        

        logic [WIDTH-1:0] out_2411;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.743)
        ) inst_2411 (
            .outp(out_2411)
        );
        

        logic [WIDTH-1:0] out_2412;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2412 (
            .a(out_3),
            .b(out_2411),
            .outp(out_2412)
        );        
        

        logic [WIDTH-1:0] out_2413;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2413 (
            .a(out_2315),
            .b(out_2412),
            .outp(out_2413)
        );        
        

        logic [WIDTH-1:0] out_2414;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.243)
        ) inst_2414 (
            .outp(out_2414)
        );
        

        logic [WIDTH-1:0] out_2415;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2415 (
            .a(out_2414),
            .b(out_3),
            .outp(out_2415)
        );        
        

        logic [WIDTH-1:0] out_2416;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2416 (
            .a(out_2413),
            .b(out_2415),
            .outp(out_2416)
        );        
        

        logic [WIDTH-1:0] out_2417;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.468)
        ) inst_2417 (
            .outp(out_2417)
        );
        

        logic [WIDTH-1:0] out_2418;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2418 (
            .a(out_3),
            .b(out_2417),
            .outp(out_2418)
        );        
        

        logic [WIDTH-1:0] out_2419;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2419 (
            .in(out_2418),
            .outp(out_2419)
        );
        

        logic [WIDTH-1:0] out_2420;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2420 (
            .a(out_753),
            .b(out_2419),
            .outp(out_2420)
        );        
        

        logic [WIDTH-1:0] out_2421;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2421 (
            .in(out_2420),
            .outp(out_2421)
        );
        

        logic [WIDTH-1:0] out_2422;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2422 (
            .a(out_2421),
            .b(out_21),
            .outp(out_2422)
        );        
        

        logic [WIDTH-1:0] out_2423;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.10808)
        ) inst_2423 (
            .outp(out_2423)
        );
        

        logic [WIDTH-1:0] out_2424;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2424 (
            .a(out_2423),
            .b(out_559),
            .outp(out_2424)
        );        
        

        logic [WIDTH-1:0] out_2425;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2425 (
            .a(out_556),
            .b(out_2424),
            .outp(out_2425)
        );        
        

        logic [WIDTH-1:0] out_2426;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2426 (
            .a(out_2290),
            .b(out_2425),
            .outp(out_2426)
        );        
        

        logic [WIDTH-1:0] out_2427;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.55693)
        ) inst_2427 (
            .outp(out_2427)
        );
        

        logic [WIDTH-1:0] out_2428;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2428 (
            .a(out_2427),
            .b(out_556),
            .outp(out_2428)
        );        
        

        logic [WIDTH-1:0] out_2429;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2429 (
            .a(out_2428),
            .b(out_566),
            .outp(out_2429)
        );        
        

        logic [WIDTH-1:0] out_2430;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2430 (
            .in(out_2429),
            .outp(out_2430)
        );
        

        logic [WIDTH-1:0] out_2431;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2431 (
            .a(out_2426),
            .b(out_2430),
            .outp(out_2431)
        );        
        

        logic [WIDTH-1:0] out_2432;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.55693)
        ) inst_2432 (
            .outp(out_2432)
        );
        

        logic [WIDTH-1:0] out_2433;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2433 (
            .a(out_2432),
            .b(out_556),
            .outp(out_2433)
        );        
        

        logic [WIDTH-1:0] out_2434;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2434 (
            .a(out_2433),
            .b(out_566),
            .outp(out_2434)
        );        
        

        logic [WIDTH-1:0] out_2435;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2435 (
            .a(out_2424),
            .b(out_556),
            .outp(out_2435)
        );        
        

        logic [WIDTH-1:0] out_2436;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2436 (
            .a(out_2434),
            .b(out_2435),
            .outp(out_2436)
        );        
        

        logic [WIDTH-1:0] out_2437;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2437 (
            .a(out_2436),
            .b(out_2300),
            .outp(out_2437)
        );        
        

        logic [WIDTH-1:0] out_2438;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2438 (
            .a(out_2431),
            .b(out_2437),
            .outp(out_2438)
        );        
        

        logic [WIDTH-1:0] out_2439;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2439 (
            .in(out_2438),
            .outp(out_2439)
        );
        

        logic [WIDTH-1:0] out_2440;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2440 (
            .a(out_2422),
            .b(out_2439),
            .outp(out_2440)
        );        
        

        logic [WIDTH-1:0] out_2441;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2441 (
            .a(out_9),
            .b(out_2421),
            .outp(out_2441)
        );        
        

        logic [WIDTH-1:0] out_2442;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2442 (
            .a(out_2440),
            .b(out_2441),
            .outp(out_2442)
        );        
        

        logic [WIDTH-1:0] out_2443;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2443 (
            .a(out_2416),
            .b(out_2442),
            .outp(out_2443)
        );        
        

        logic [WIDTH-1:0] out_2444;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2444 (
            .a(out_2422),
            .b(out_2443),
            .outp(out_2444)
        );        
        

        logic [WIDTH-1:0] out_2445;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2445 (
            .a(out_2410),
            .b(out_2444),
            .outp(out_2445)
        );        
        

        logic [WIDTH-1:0] out_2446;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.475)
        ) inst_2446 (
            .outp(out_2446)
        );
        

        logic [WIDTH-1:0] out_2447;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2447 (
            .a(out_2446),
            .b(out_14),
            .outp(out_2447)
        );        
        

        logic [WIDTH-1:0] out_2448;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2448 (
            .in(out_2447),
            .outp(out_2448)
        );
        

        logic [WIDTH-1:0] out_2449;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2449 (
            .a(out_727),
            .b(out_2448),
            .outp(out_2449)
        );        
        

        logic [WIDTH-1:0] out_2450;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.643001)
        ) inst_2450 (
            .outp(out_2450)
        );
        

        logic [WIDTH-1:0] out_2451;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2451 (
            .a(out_3),
            .b(out_2450),
            .outp(out_2451)
        );        
        

        logic [WIDTH-1:0] out_2452;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2452 (
            .a(out_2449),
            .b(out_2451),
            .outp(out_2452)
        );        
        

        logic [WIDTH-1:0] out_2453;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.543)
        ) inst_2453 (
            .outp(out_2453)
        );
        

        logic [WIDTH-1:0] out_2454;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2454 (
            .a(out_2453),
            .b(out_3),
            .outp(out_2454)
        );        
        

        logic [WIDTH-1:0] out_2455;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2455 (
            .a(out_2452),
            .b(out_2454),
            .outp(out_2455)
        );        
        

        logic [WIDTH-1:0] out_2456;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2456 (
            .a(out_2445),
            .b(out_2455),
            .outp(out_2456)
        );        
        

        logic [WIDTH-1:0] out_2457;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.818)
        ) inst_2457 (
            .outp(out_2457)
        );
        

        logic [WIDTH-1:0] out_2458;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2458 (
            .a(out_3),
            .b(out_2457),
            .outp(out_2458)
        );        
        

        logic [WIDTH-1:0] out_2459;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2459 (
            .in(out_2458),
            .outp(out_2459)
        );
        

        logic [WIDTH-1:0] out_2460;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2460 (
            .a(out_753),
            .b(out_2459),
            .outp(out_2460)
        );        
        

        logic [WIDTH-1:0] out_2461;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2461 (
            .in(out_2460),
            .outp(out_2461)
        );
        

        logic [WIDTH-1:0] out_2462;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2462 (
            .a(out_9),
            .b(out_2461),
            .outp(out_2462)
        );        
        

        logic [WIDTH-1:0] out_2463;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2463 (
            .a(out_2461),
            .b(out_21),
            .outp(out_2463)
        );        
        

        logic [WIDTH-1:0] out_2464;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2464 (
            .a(out_2462),
            .b(out_2463),
            .outp(out_2464)
        );        
        

        logic [WIDTH-1:0] out_2465;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2465 (
            .a(out_2456),
            .b(out_2464),
            .outp(out_2465)
        );        
        

        logic [WIDTH-1:0] out_2466;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.937)
        ) inst_2466 (
            .outp(out_2466)
        );
        

        logic [WIDTH-1:0] out_2467;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2467 (
            .a(out_2466),
            .b(out_3),
            .outp(out_2467)
        );        
        

        logic [WIDTH-1:0] out_2468;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2468 (
            .in(out_2467),
            .outp(out_2468)
        );
        

        logic [WIDTH-1:0] out_2469;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.34167)
        ) inst_2469 (
            .outp(out_2469)
        );
        

        logic [WIDTH-1:0] out_2470;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2470 (
            .a(out_2469),
            .b(out_1933),
            .outp(out_2470)
        );        
        

        logic [WIDTH-1:0] out_2471;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2471 (
            .in(out_2470),
            .outp(out_2471)
        );
        

        logic [WIDTH-1:0] out_2472;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2472 (
            .a(out_2468),
            .b(out_2471),
            .outp(out_2472)
        );        
        

        logic [WIDTH-1:0] out_2473;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2473 (
            .in(out_2472),
            .outp(out_2473)
        );
        

        logic [WIDTH-1:0] out_2474;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2474 (
            .a(out_2473),
            .b(out_460),
            .outp(out_2474)
        );        
        

        logic [WIDTH-1:0] out_2475;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.3292)
        ) inst_2475 (
            .outp(out_2475)
        );
        

        logic [WIDTH-1:0] out_2476;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2476 (
            .a(out_2475),
            .b(out_1891),
            .outp(out_2476)
        );        
        

        logic [WIDTH-1:0] out_2477;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2477 (
            .a(out_2476),
            .b(out_137),
            .outp(out_2477)
        );        
        

        logic [WIDTH-1:0] out_2478;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2527)
        ) inst_2478 (
            .outp(out_2478)
        );
        

        logic [WIDTH-1:0] out_2479;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2479 (
            .a(out_1897),
            .b(out_2478),
            .outp(out_2479)
        );        
        

        logic [WIDTH-1:0] out_2480;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2480 (
            .a(out_2479),
            .b(out_566),
            .outp(out_2480)
        );        
        

        logic [WIDTH-1:0] out_2481;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2481 (
            .in(out_2480),
            .outp(out_2481)
        );
        

        logic [WIDTH-1:0] out_2482;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2482 (
            .a(out_2477),
            .b(out_2481),
            .outp(out_2482)
        );        
        

        logic [WIDTH-1:0] out_2483;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.726)
        ) inst_2483 (
            .outp(out_2483)
        );
        

        logic [WIDTH-1:0] out_2484;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2484 (
            .a(out_2483),
            .b(out_1904),
            .outp(out_2484)
        );        
        

        logic [WIDTH-1:0] out_2485;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2485 (
            .a(out_2484),
            .b(out_1907),
            .outp(out_2485)
        );        
        

        logic [WIDTH-1:0] out_2486;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2486 (
            .a(out_2482),
            .b(out_2485),
            .outp(out_2486)
        );        
        

        logic [WIDTH-1:0] out_2487;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2487 (
            .a(out_1907),
            .b(out_2484),
            .outp(out_2487)
        );        
        

        logic [WIDTH-1:0] out_2488;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2527)
        ) inst_2488 (
            .outp(out_2488)
        );
        

        logic [WIDTH-1:0] out_2489;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2489 (
            .a(out_1897),
            .b(out_2488),
            .outp(out_2489)
        );        
        

        logic [WIDTH-1:0] out_2490;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2490 (
            .a(out_2489),
            .b(out_566),
            .outp(out_2490)
        );        
        

        logic [WIDTH-1:0] out_2491;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2491 (
            .a(out_2487),
            .b(out_2490),
            .outp(out_2491)
        );        
        

        logic [WIDTH-1:0] out_2492;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2492 (
            .a(out_137),
            .b(out_2476),
            .outp(out_2492)
        );        
        

        logic [WIDTH-1:0] out_2493;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2493 (
            .a(out_2491),
            .b(out_2492),
            .outp(out_2493)
        );        
        

        logic [WIDTH-1:0] out_2494;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2494 (
            .a(out_2486),
            .b(out_2493),
            .outp(out_2494)
        );        
        

        logic [WIDTH-1:0] out_2495;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2495 (
            .in(out_2494),
            .outp(out_2495)
        );
        

        logic [WIDTH-1:0] out_2496;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2496 (
            .a(out_2474),
            .b(out_2495),
            .outp(out_2496)
        );        
        

        logic [WIDTH-1:0] out_2497;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2497 (
            .a(out_31),
            .b(out_14),
            .outp(out_2497)
        );        
        

        logic [WIDTH-1:0] out_2498;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2498 (
            .a(out_2496),
            .b(out_2497),
            .outp(out_2498)
        );        
        

        logic [WIDTH-1:0] out_2499;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.25)
        ) inst_2499 (
            .outp(out_2499)
        );
        

        logic [WIDTH-1:0] out_2500;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2500 (
            .a(out_2499),
            .b(out_14),
            .outp(out_2500)
        );        
        

        logic [WIDTH-1:0] out_2501;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2501 (
            .in(out_2500),
            .outp(out_2501)
        );
        

        logic [WIDTH-1:0] out_2502;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2502 (
            .a(out_2498),
            .b(out_2501),
            .outp(out_2502)
        );        
        

        logic [WIDTH-1:0] out_2503;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.862)
        ) inst_2503 (
            .outp(out_2503)
        );
        

        logic [WIDTH-1:0] out_2504;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2504 (
            .a(out_2503),
            .b(out_3),
            .outp(out_2504)
        );        
        

        logic [WIDTH-1:0] out_2505;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2505 (
            .a(out_2502),
            .b(out_2504),
            .outp(out_2505)
        );        
        

        logic [WIDTH-1:0] out_2506;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.012)
        ) inst_2506 (
            .outp(out_2506)
        );
        

        logic [WIDTH-1:0] out_2507;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2507 (
            .a(out_2506),
            .b(out_3),
            .outp(out_2507)
        );        
        

        logic [WIDTH-1:0] out_2508;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2508 (
            .in(out_2507),
            .outp(out_2508)
        );
        

        logic [WIDTH-1:0] out_2509;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2509 (
            .a(out_2505),
            .b(out_2508),
            .outp(out_2509)
        );        
        

        logic [WIDTH-1:0] out_2510;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2510 (
            .a(out_2465),
            .b(out_2509),
            .outp(out_2510)
        );        
        

        logic [WIDTH-1:0] out_2511;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2511 (
            .in(out_2497),
            .outp(out_2511)
        );
        

        logic [WIDTH-1:0] out_2512;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.912)
        ) inst_2512 (
            .outp(out_2512)
        );
        

        logic [WIDTH-1:0] out_2513;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2513 (
            .a(out_2512),
            .b(out_3),
            .outp(out_2513)
        );        
        

        logic [WIDTH-1:0] out_2514;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2514 (
            .in(out_2513),
            .outp(out_2514)
        );
        

        logic [WIDTH-1:0] out_2515;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2515 (
            .a(out_2511),
            .b(out_2514),
            .outp(out_2515)
        );        
        

        logic [WIDTH-1:0] out_2516;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2516 (
            .in(out_2515),
            .outp(out_2516)
        );
        

        logic [WIDTH-1:0] out_2517;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2517 (
            .a(out_2516),
            .b(out_460),
            .outp(out_2517)
        );        
        

        logic [WIDTH-1:0] out_2518;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2518 (
            .a(out_2510),
            .b(out_2517),
            .outp(out_2518)
        );        
        

        logic [WIDTH-1:0] out_2519;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.162)
        ) inst_2519 (
            .outp(out_2519)
        );
        

        logic [WIDTH-1:0] out_2520;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2520 (
            .a(out_2519),
            .b(out_3),
            .outp(out_2520)
        );        
        

        logic [WIDTH-1:0] out_2521;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2521 (
            .a(out_2094),
            .b(out_2520),
            .outp(out_2521)
        );        
        

        logic [WIDTH-1:0] out_2522;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.262)
        ) inst_2522 (
            .outp(out_2522)
        );
        

        logic [WIDTH-1:0] out_2523;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2523 (
            .a(out_2522),
            .b(out_3),
            .outp(out_2523)
        );        
        

        logic [WIDTH-1:0] out_2524;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2524 (
            .in(out_2523),
            .outp(out_2524)
        );
        

        logic [WIDTH-1:0] out_2525;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2525 (
            .a(out_2521),
            .b(out_2524),
            .outp(out_2525)
        );        
        

        logic [WIDTH-1:0] out_2526;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2526 (
            .a(out_2518),
            .b(out_2525),
            .outp(out_2526)
        );        
        

        logic [WIDTH-1:0] out_2527;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.612)
        ) inst_2527 (
            .outp(out_2527)
        );
        

        logic [WIDTH-1:0] out_2528;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2528 (
            .a(out_2527),
            .b(out_3),
            .outp(out_2528)
        );        
        

        logic [WIDTH-1:0] out_2529;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2529 (
            .a(out_718),
            .b(out_2528),
            .outp(out_2529)
        );        
        

        logic [WIDTH-1:0] out_2530;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.712)
        ) inst_2530 (
            .outp(out_2530)
        );
        

        logic [WIDTH-1:0] out_2531;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2531 (
            .a(out_2530),
            .b(out_3),
            .outp(out_2531)
        );        
        

        logic [WIDTH-1:0] out_2532;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2532 (
            .in(out_2531),
            .outp(out_2532)
        );
        

        logic [WIDTH-1:0] out_2533;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2533 (
            .a(out_2529),
            .b(out_2532),
            .outp(out_2533)
        );        
        

        logic [WIDTH-1:0] out_2534;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2534 (
            .a(out_2526),
            .b(out_2533),
            .outp(out_2534)
        );        
        

        logic [WIDTH-1:0] out_2535;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2535 (
            .a(out_727),
            .b(out_2113),
            .outp(out_2535)
        );        
        

        logic [WIDTH-1:0] out_2536;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2536 (
            .a(out_2535),
            .b(out_2520),
            .outp(out_2536)
        );        
        

        logic [WIDTH-1:0] out_2537;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2537 (
            .a(out_2536),
            .b(out_2532),
            .outp(out_2537)
        );        
        

        logic [WIDTH-1:0] out_2538;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.437)
        ) inst_2538 (
            .outp(out_2538)
        );
        

        logic [WIDTH-1:0] out_2539;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2539 (
            .a(out_2538),
            .b(out_3),
            .outp(out_2539)
        );        
        

        logic [WIDTH-1:0] out_2540;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2540 (
            .in(out_2539),
            .outp(out_2540)
        );
        

        logic [WIDTH-1:0] out_2541;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2541 (
            .a(out_753),
            .b(out_2540),
            .outp(out_2541)
        );        
        

        logic [WIDTH-1:0] out_2542;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2542 (
            .in(out_2541),
            .outp(out_2542)
        );
        

        logic [WIDTH-1:0] out_2543;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2543 (
            .a(out_9),
            .b(out_2542),
            .outp(out_2543)
        );        
        

        logic [WIDTH-1:0] out_2544;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2544 (
            .a(out_2537),
            .b(out_2543),
            .outp(out_2544)
        );        
        

        logic [WIDTH-1:0] out_2545;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2545 (
            .a(out_2542),
            .b(out_21),
            .outp(out_2545)
        );        
        

        logic [WIDTH-1:0] out_2546;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2546 (
            .a(out_2544),
            .b(out_2545),
            .outp(out_2546)
        );        
        

        logic [WIDTH-1:0] out_2547;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2547 (
            .a(out_2534),
            .b(out_2546),
            .outp(out_2547)
        );        
        

        logic [WIDTH-1:0] out_2548;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.962)
        ) inst_2548 (
            .outp(out_2548)
        );
        

        logic [WIDTH-1:0] out_2549;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2549 (
            .a(out_2548),
            .b(out_3),
            .outp(out_2549)
        );        
        

        logic [WIDTH-1:0] out_2550;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2550 (
            .a(out_2128),
            .b(out_2549),
            .outp(out_2550)
        );        
        

        logic [WIDTH-1:0] out_2551;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.062)
        ) inst_2551 (
            .outp(out_2551)
        );
        

        logic [WIDTH-1:0] out_2552;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2552 (
            .a(out_2551),
            .b(out_3),
            .outp(out_2552)
        );        
        

        logic [WIDTH-1:0] out_2553;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2553 (
            .in(out_2552),
            .outp(out_2553)
        );
        

        logic [WIDTH-1:0] out_2554;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2554 (
            .a(out_2550),
            .b(out_2553),
            .outp(out_2554)
        );        
        

        logic [WIDTH-1:0] out_2555;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2555 (
            .a(out_2547),
            .b(out_2554),
            .outp(out_2555)
        );        
        

        logic [WIDTH-1:0] out_2556;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.812)
        ) inst_2556 (
            .outp(out_2556)
        );
        

        logic [WIDTH-1:0] out_2557;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2557 (
            .a(out_2556),
            .b(out_3),
            .outp(out_2557)
        );        
        

        logic [WIDTH-1:0] out_2558;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2558 (
            .a(out_2141),
            .b(out_2557),
            .outp(out_2558)
        );        
        

        logic [WIDTH-1:0] out_2559;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.212)
        ) inst_2559 (
            .outp(out_2559)
        );
        

        logic [WIDTH-1:0] out_2560;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2560 (
            .a(out_2559),
            .b(out_3),
            .outp(out_2560)
        );        
        

        logic [WIDTH-1:0] out_2561;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2561 (
            .in(out_2560),
            .outp(out_2561)
        );
        

        logic [WIDTH-1:0] out_2562;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2562 (
            .a(out_2558),
            .b(out_2561),
            .outp(out_2562)
        );        
        

        logic [WIDTH-1:0] out_2563;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2563 (
            .a(out_2555),
            .b(out_2562),
            .outp(out_2563)
        );        
        

        logic [WIDTH-1:0] out_2564;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2564 (
            .a(out_2149),
            .b(out_2557),
            .outp(out_2564)
        );        
        

        logic [WIDTH-1:0] out_2565;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2565 (
            .a(out_2564),
            .b(out_2561),
            .outp(out_2565)
        );        
        

        logic [WIDTH-1:0] out_2566;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2566 (
            .in(out_2557),
            .outp(out_2566)
        );
        

        logic [WIDTH-1:0] out_2567;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2567 (
            .a(out_2152),
            .b(out_2566),
            .outp(out_2567)
        );        
        

        logic [WIDTH-1:0] out_2568;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2568 (
            .in(out_2567),
            .outp(out_2568)
        );
        

        logic [WIDTH-1:0] out_2569;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2569 (
            .a(out_336),
            .b(out_2568),
            .outp(out_2569)
        );        
        

        logic [WIDTH-1:0] out_2570;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2570 (
            .a(out_2565),
            .b(out_2569),
            .outp(out_2570)
        );        
        

        logic [WIDTH-1:0] out_2571;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2571 (
            .a(out_2568),
            .b(out_343),
            .outp(out_2571)
        );        
        

        logic [WIDTH-1:0] out_2572;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2572 (
            .a(out_2570),
            .b(out_2571),
            .outp(out_2572)
        );        
        

        logic [WIDTH-1:0] out_2573;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2573 (
            .a(out_2563),
            .b(out_2572),
            .outp(out_2573)
        );        
        

        logic [WIDTH-1:0] out_2574;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.57)
        ) inst_2574 (
            .outp(out_2574)
        );
        

        logic [WIDTH-1:0] out_2575;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2575 (
            .a(out_2574),
            .b(out_3),
            .outp(out_2575)
        );        
        

        logic [WIDTH-1:0] out_2576;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2576 (
            .a(out_2161),
            .b(out_2575),
            .outp(out_2576)
        );        
        

        logic [WIDTH-1:0] out_2577;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.67)
        ) inst_2577 (
            .outp(out_2577)
        );
        

        logic [WIDTH-1:0] out_2578;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2578 (
            .a(out_2577),
            .b(out_3),
            .outp(out_2578)
        );        
        

        logic [WIDTH-1:0] out_2579;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2579 (
            .in(out_2578),
            .outp(out_2579)
        );
        

        logic [WIDTH-1:0] out_2580;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2580 (
            .a(out_2576),
            .b(out_2579),
            .outp(out_2580)
        );        
        

        logic [WIDTH-1:0] out_2581;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2581 (
            .a(out_2573),
            .b(out_2580),
            .outp(out_2581)
        );        
        

        logic [WIDTH-1:0] out_2582;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2582 (
            .a(out_718),
            .b(out_2404),
            .outp(out_2582)
        );        
        

        logic [WIDTH-1:0] out_2583;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.182)
        ) inst_2583 (
            .outp(out_2583)
        );
        

        logic [WIDTH-1:0] out_2584;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2584 (
            .a(out_2583),
            .b(out_3),
            .outp(out_2584)
        );        
        

        logic [WIDTH-1:0] out_2585;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2585 (
            .in(out_2584),
            .outp(out_2585)
        );
        

        logic [WIDTH-1:0] out_2586;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2586 (
            .a(out_2582),
            .b(out_2585),
            .outp(out_2586)
        );        
        

        logic [WIDTH-1:0] out_2587;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2587 (
            .in(out_2405),
            .outp(out_2587)
        );
        

        logic [WIDTH-1:0] out_2588;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2588 (
            .a(out_753),
            .b(out_2587),
            .outp(out_2588)
        );        
        

        logic [WIDTH-1:0] out_2589;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2589 (
            .in(out_2588),
            .outp(out_2589)
        );
        

        logic [WIDTH-1:0] out_2590;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2590 (
            .a(out_9),
            .b(out_2589),
            .outp(out_2590)
        );        
        

        logic [WIDTH-1:0] out_2591;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2591 (
            .a(out_2586),
            .b(out_2590),
            .outp(out_2591)
        );        
        

        logic [WIDTH-1:0] out_2592;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2592 (
            .a(out_2589),
            .b(out_21),
            .outp(out_2592)
        );        
        

        logic [WIDTH-1:0] out_2593;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2593 (
            .a(out_2591),
            .b(out_2592),
            .outp(out_2593)
        );        
        

        logic [WIDTH-1:0] out_2594;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2594 (
            .a(out_2581),
            .b(out_2593),
            .outp(out_2594)
        );        
        

        logic [WIDTH-1:0] out_2595;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.807)
        ) inst_2595 (
            .outp(out_2595)
        );
        

        logic [WIDTH-1:0] out_2596;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2596 (
            .a(out_2595),
            .b(out_3),
            .outp(out_2596)
        );        
        

        logic [WIDTH-1:0] out_2597;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2597 (
            .a(out_2240),
            .b(out_2596),
            .outp(out_2597)
        );        
        

        logic [WIDTH-1:0] out_2598;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.907)
        ) inst_2598 (
            .outp(out_2598)
        );
        

        logic [WIDTH-1:0] out_2599;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2599 (
            .a(out_2598),
            .b(out_3),
            .outp(out_2599)
        );        
        

        logic [WIDTH-1:0] out_2600;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2600 (
            .in(out_2599),
            .outp(out_2600)
        );
        

        logic [WIDTH-1:0] out_2601;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2601 (
            .a(out_2597),
            .b(out_2600),
            .outp(out_2601)
        );        
        

        logic [WIDTH-1:0] out_2602;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2602 (
            .a(out_2594),
            .b(out_2601),
            .outp(out_2602)
        );        
        

        logic [WIDTH-1:0] out_2603;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.257)
        ) inst_2603 (
            .outp(out_2603)
        );
        

        logic [WIDTH-1:0] out_2604;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2604 (
            .a(out_2603),
            .b(out_3),
            .outp(out_2604)
        );        
        

        logic [WIDTH-1:0] out_2605;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2605 (
            .a(out_2161),
            .b(out_2604),
            .outp(out_2605)
        );        
        

        logic [WIDTH-1:0] out_2606;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.357)
        ) inst_2606 (
            .outp(out_2606)
        );
        

        logic [WIDTH-1:0] out_2607;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2607 (
            .a(out_2606),
            .b(out_3),
            .outp(out_2607)
        );        
        

        logic [WIDTH-1:0] out_2608;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2608 (
            .in(out_2607),
            .outp(out_2608)
        );
        

        logic [WIDTH-1:0] out_2609;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2609 (
            .a(out_2605),
            .b(out_2608),
            .outp(out_2609)
        );        
        

        logic [WIDTH-1:0] out_2610;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2610 (
            .a(out_2602),
            .b(out_2609),
            .outp(out_2610)
        );        
        

        logic [WIDTH-1:0] out_2611;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2611 (
            .a(out_727),
            .b(out_2259),
            .outp(out_2611)
        );        
        

        logic [WIDTH-1:0] out_2612;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2612 (
            .a(out_2611),
            .b(out_2596),
            .outp(out_2612)
        );        
        

        logic [WIDTH-1:0] out_2613;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2613 (
            .a(out_2612),
            .b(out_2608),
            .outp(out_2613)
        );        
        

        logic [WIDTH-1:0] out_2614;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.082)
        ) inst_2614 (
            .outp(out_2614)
        );
        

        logic [WIDTH-1:0] out_2615;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2615 (
            .a(out_2614),
            .b(out_3),
            .outp(out_2615)
        );        
        

        logic [WIDTH-1:0] out_2616;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2616 (
            .in(out_2615),
            .outp(out_2616)
        );
        

        logic [WIDTH-1:0] out_2617;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2617 (
            .a(out_753),
            .b(out_2616),
            .outp(out_2617)
        );        
        

        logic [WIDTH-1:0] out_2618;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2618 (
            .in(out_2617),
            .outp(out_2618)
        );
        

        logic [WIDTH-1:0] out_2619;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2619 (
            .a(out_9),
            .b(out_2618),
            .outp(out_2619)
        );        
        

        logic [WIDTH-1:0] out_2620;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2620 (
            .a(out_2613),
            .b(out_2619),
            .outp(out_2620)
        );        
        

        logic [WIDTH-1:0] out_2621;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2621 (
            .a(out_2618),
            .b(out_21),
            .outp(out_2621)
        );        
        

        logic [WIDTH-1:0] out_2622;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2622 (
            .a(out_2620),
            .b(out_2621),
            .outp(out_2622)
        );        
        

        logic [WIDTH-1:0] out_2623;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2623 (
            .a(out_2610),
            .b(out_2622),
            .outp(out_2623)
        );        
        

        logic [WIDTH-1:0] out_2624;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.477)
        ) inst_2624 (
            .outp(out_2624)
        );
        

        logic [WIDTH-1:0] out_2625;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2625 (
            .a(out_2624),
            .b(out_3),
            .outp(out_2625)
        );        
        

        logic [WIDTH-1:0] out_2626;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2626 (
            .a(out_2273),
            .b(out_2625),
            .outp(out_2626)
        );        
        

        logic [WIDTH-1:0] out_2627;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.577)
        ) inst_2627 (
            .outp(out_2627)
        );
        

        logic [WIDTH-1:0] out_2628;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2628 (
            .a(out_2627),
            .b(out_3),
            .outp(out_2628)
        );        
        

        logic [WIDTH-1:0] out_2629;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2629 (
            .in(out_2628),
            .outp(out_2629)
        );
        

        logic [WIDTH-1:0] out_2630;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2630 (
            .a(out_2626),
            .b(out_2629),
            .outp(out_2630)
        );        
        

        logic [WIDTH-1:0] out_2631;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2631 (
            .a(out_2623),
            .b(out_2630),
            .outp(out_2631)
        );        
        

        logic [WIDTH-1:0] out_2632;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.66557)
        ) inst_2632 (
            .outp(out_2632)
        );
        

        logic [WIDTH-1:0] out_2633;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2633 (
            .a(out_2632),
            .b(out_3),
            .outp(out_2633)
        );        
        

        logic [WIDTH-1:0] out_2634;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2634 (
            .a(out_2633),
            .b(out_1495),
            .outp(out_2634)
        );        
        

        logic [WIDTH-1:0] out_2635;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2635 (
            .in(out_2634),
            .outp(out_2635)
        );
        

        logic [WIDTH-1:0] out_2636;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2636 (
            .a(out_753),
            .b(out_2635),
            .outp(out_2636)
        );        
        

        logic [WIDTH-1:0] out_2637;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2637 (
            .in(out_2636),
            .outp(out_2637)
        );
        

        logic [WIDTH-1:0] out_2638;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2638 (
            .a(out_9),
            .b(out_2637),
            .outp(out_2638)
        );        
        

        logic [WIDTH-1:0] out_2639;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2639 (
            .a(out_2637),
            .b(out_21),
            .outp(out_2639)
        );        
        

        logic [WIDTH-1:0] out_2640;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2640 (
            .a(out_2638),
            .b(out_2639),
            .outp(out_2640)
        );        
        

        logic [WIDTH-1:0] out_2641;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2641 (
            .a(out_2631),
            .b(out_2640),
            .outp(out_2641)
        );        
        

        logic [WIDTH-1:0] out_2642;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.9605)
        ) inst_2642 (
            .outp(out_2642)
        );
        

        logic [WIDTH-1:0] out_2643;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2643 (
            .a(out_3),
            .b(out_2642),
            .outp(out_2643)
        );        
        

        logic [WIDTH-1:0] out_2644;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2644 (
            .in(out_2643),
            .outp(out_2644)
        );
        

        logic [WIDTH-1:0] out_2645;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2645 (
            .a(out_1300),
            .b(out_2644),
            .outp(out_2645)
        );        
        

        logic [WIDTH-1:0] out_2646;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2646 (
            .in(out_2645),
            .outp(out_2646)
        );
        

        logic [WIDTH-1:0] out_2647;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2647 (
            .a(out_2646),
            .b(out_21),
            .outp(out_2647)
        );        
        

        logic [WIDTH-1:0] out_2648;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.17851)
        ) inst_2648 (
            .outp(out_2648)
        );
        

        logic [WIDTH-1:0] out_2649;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2649 (
            .a(out_559),
            .b(out_2648),
            .outp(out_2649)
        );        
        

        logic [WIDTH-1:0] out_2650;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2650 (
            .a(out_556),
            .b(out_2649),
            .outp(out_2650)
        );        
        

        logic [WIDTH-1:0] out_2651;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2651 (
            .a(out_1806),
            .b(out_2650),
            .outp(out_2651)
        );        
        

        logic [WIDTH-1:0] out_2652;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.228514)
        ) inst_2652 (
            .outp(out_2652)
        );
        

        logic [WIDTH-1:0] out_2653;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2653 (
            .a(out_556),
            .b(out_566),
            .outp(out_2653)
        );        
        

        logic [WIDTH-1:0] out_2654;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2654 (
            .a(out_2652),
            .b(out_2653),
            .outp(out_2654)
        );        
        

        logic [WIDTH-1:0] out_2655;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2655 (
            .a(out_2651),
            .b(out_2654),
            .outp(out_2655)
        );        
        

        logic [WIDTH-1:0] out_2656;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2656 (
            .a(out_2653),
            .b(out_2652),
            .outp(out_2656)
        );        
        

        logic [WIDTH-1:0] out_2657;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2657 (
            .a(out_2649),
            .b(out_556),
            .outp(out_2657)
        );        
        

        logic [WIDTH-1:0] out_2658;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2658 (
            .a(out_2656),
            .b(out_2657),
            .outp(out_2658)
        );        
        

        logic [WIDTH-1:0] out_2659;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2659 (
            .a(out_2658),
            .b(out_1813),
            .outp(out_2659)
        );        
        

        logic [WIDTH-1:0] out_2660;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2660 (
            .a(out_2655),
            .b(out_2659),
            .outp(out_2660)
        );        
        

        logic [WIDTH-1:0] out_2661;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2661 (
            .in(out_2660),
            .outp(out_2661)
        );
        

        logic [WIDTH-1:0] out_2662;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2662 (
            .a(out_2647),
            .b(out_2661),
            .outp(out_2662)
        );        
        

        logic [WIDTH-1:0] out_2663;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2663 (
            .a(out_9),
            .b(out_2646),
            .outp(out_2663)
        );        
        

        logic [WIDTH-1:0] out_2664;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2664 (
            .a(out_2662),
            .b(out_2663),
            .outp(out_2664)
        );        
        

        logic [WIDTH-1:0] out_2665;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2665 (
            .a(out_1785),
            .b(out_1789),
            .outp(out_2665)
        );        
        

        logic [WIDTH-1:0] out_2666;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.23551)
        ) inst_2666 (
            .outp(out_2666)
        );
        

        logic [WIDTH-1:0] out_2667;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2667 (
            .a(out_3),
            .b(out_2666),
            .outp(out_2667)
        );        
        

        logic [WIDTH-1:0] out_2668;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2668 (
            .a(out_2665),
            .b(out_2667),
            .outp(out_2668)
        );        
        

        logic [WIDTH-1:0] out_2669;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.73551)
        ) inst_2669 (
            .outp(out_2669)
        );
        

        logic [WIDTH-1:0] out_2670;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2670 (
            .a(out_2669),
            .b(out_3),
            .outp(out_2670)
        );        
        

        logic [WIDTH-1:0] out_2671;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2671 (
            .a(out_2668),
            .b(out_2670),
            .outp(out_2671)
        );        
        

        logic [WIDTH-1:0] out_2672;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2672 (
            .a(out_2664),
            .b(out_2671),
            .outp(out_2672)
        );        
        

        logic [WIDTH-1:0] out_2673;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2673 (
            .a(out_2672),
            .b(out_2647),
            .outp(out_2673)
        );        
        

        logic [WIDTH-1:0] out_2674;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2674 (
            .a(out_2641),
            .b(out_2673),
            .outp(out_2674)
        );        
        

        logic [WIDTH-1:0] out_2675;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.5355)
        ) inst_2675 (
            .outp(out_2675)
        );
        

        logic [WIDTH-1:0] out_2676;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2676 (
            .a(out_3),
            .b(out_2675),
            .outp(out_2676)
        );        
        

        logic [WIDTH-1:0] out_2677;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2677 (
            .a(out_1244),
            .b(out_2676),
            .outp(out_2677)
        );        
        

        logic [WIDTH-1:0] out_2678;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.4355)
        ) inst_2678 (
            .outp(out_2678)
        );
        

        logic [WIDTH-1:0] out_2679;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2679 (
            .a(out_2678),
            .b(out_3),
            .outp(out_2679)
        );        
        

        logic [WIDTH-1:0] out_2680;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2680 (
            .a(out_2677),
            .b(out_2679),
            .outp(out_2680)
        );        
        

        logic [WIDTH-1:0] out_2681;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2681 (
            .a(out_2680),
            .b(out_1299),
            .outp(out_2681)
        );        
        

        logic [WIDTH-1:0] out_2682;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2682 (
            .a(out_2674),
            .b(out_2681),
            .outp(out_2682)
        );        
        

        logic [WIDTH-1:0] out_2683;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2683 (
            .a(out_1244),
            .b(out_1324),
            .outp(out_2683)
        );        
        

        logic [WIDTH-1:0] out_2684;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.0855)
        ) inst_2684 (
            .outp(out_2684)
        );
        

        logic [WIDTH-1:0] out_2685;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2685 (
            .a(out_3),
            .b(out_2684),
            .outp(out_2685)
        );        
        

        logic [WIDTH-1:0] out_2686;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2686 (
            .a(out_2683),
            .b(out_2685),
            .outp(out_2686)
        );        
        

        logic [WIDTH-1:0] out_2687;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.9855)
        ) inst_2687 (
            .outp(out_2687)
        );
        

        logic [WIDTH-1:0] out_2688;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2688 (
            .a(out_2687),
            .b(out_3),
            .outp(out_2688)
        );        
        

        logic [WIDTH-1:0] out_2689;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2689 (
            .a(out_2686),
            .b(out_2688),
            .outp(out_2689)
        );        
        

        logic [WIDTH-1:0] out_2690;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2690 (
            .a(out_2682),
            .b(out_2689),
            .outp(out_2690)
        );        
        

        logic [WIDTH-1:0] out_2691;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2691 (
            .a(out_2676),
            .b(out_2688),
            .outp(out_2691)
        );        
        

        logic [WIDTH-1:0] out_2692;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2692 (
            .a(out_2691),
            .b(out_1338),
            .outp(out_2692)
        );        
        

        logic [WIDTH-1:0] out_2693;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2693 (
            .a(out_2692),
            .b(out_1342),
            .outp(out_2693)
        );        
        

        logic [WIDTH-1:0] out_2694;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.2605)
        ) inst_2694 (
            .outp(out_2694)
        );
        

        logic [WIDTH-1:0] out_2695;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2695 (
            .a(out_3),
            .b(out_2694),
            .outp(out_2695)
        );        
        

        logic [WIDTH-1:0] out_2696;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2696 (
            .in(out_2695),
            .outp(out_2696)
        );
        

        logic [WIDTH-1:0] out_2697;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2697 (
            .a(out_2696),
            .b(out_1300),
            .outp(out_2697)
        );        
        

        logic [WIDTH-1:0] out_2698;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2698 (
            .in(out_2697),
            .outp(out_2698)
        );
        

        logic [WIDTH-1:0] out_2699;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2699 (
            .a(out_9),
            .b(out_2698),
            .outp(out_2699)
        );        
        

        logic [WIDTH-1:0] out_2700;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2700 (
            .a(out_2693),
            .b(out_2699),
            .outp(out_2700)
        );        
        

        logic [WIDTH-1:0] out_2701;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2701 (
            .a(out_2698),
            .b(out_21),
            .outp(out_2701)
        );        
        

        logic [WIDTH-1:0] out_2702;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2702 (
            .a(out_2700),
            .b(out_2701),
            .outp(out_2702)
        );        
        

        logic [WIDTH-1:0] out_2703;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2703 (
            .a(out_2690),
            .b(out_2702),
            .outp(out_2703)
        );        
        

        logic [WIDTH-1:0] out_2704;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2704 (
            .a(out_1324),
            .b(out_1513),
            .outp(out_2704)
        );        
        

        logic [WIDTH-1:0] out_2705;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.7355)
        ) inst_2705 (
            .outp(out_2705)
        );
        

        logic [WIDTH-1:0] out_2706;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2706 (
            .a(out_3),
            .b(out_2705),
            .outp(out_2706)
        );        
        

        logic [WIDTH-1:0] out_2707;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2707 (
            .a(out_2704),
            .b(out_2706),
            .outp(out_2707)
        );        
        

        logic [WIDTH-1:0] out_2708;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.6355)
        ) inst_2708 (
            .outp(out_2708)
        );
        

        logic [WIDTH-1:0] out_2709;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2709 (
            .a(out_2708),
            .b(out_3),
            .outp(out_2709)
        );        
        

        logic [WIDTH-1:0] out_2710;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2710 (
            .a(out_2707),
            .b(out_2709),
            .outp(out_2710)
        );        
        

        logic [WIDTH-1:0] out_2711;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2711 (
            .a(out_2703),
            .b(out_2710),
            .outp(out_2711)
        );        
        

        logic [WIDTH-1:0] out_2712;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2712 (
            .a(out_1292),
            .b(out_1525),
            .outp(out_2712)
        );        
        

        logic [WIDTH-1:0] out_2713;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.8855)
        ) inst_2713 (
            .outp(out_2713)
        );
        

        logic [WIDTH-1:0] out_2714;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2714 (
            .a(out_3),
            .b(out_2713),
            .outp(out_2714)
        );        
        

        logic [WIDTH-1:0] out_2715;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2715 (
            .a(out_2712),
            .b(out_2714),
            .outp(out_2715)
        );        
        

        logic [WIDTH-1:0] out_2716;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.4855)
        ) inst_2716 (
            .outp(out_2716)
        );
        

        logic [WIDTH-1:0] out_2717;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2717 (
            .a(out_2716),
            .b(out_3),
            .outp(out_2717)
        );        
        

        logic [WIDTH-1:0] out_2718;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2718 (
            .a(out_2715),
            .b(out_2717),
            .outp(out_2718)
        );        
        

        logic [WIDTH-1:0] out_2719;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2719 (
            .a(out_2711),
            .b(out_2718),
            .outp(out_2719)
        );        
        

        logic [WIDTH-1:0] out_2720;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2720 (
            .a(out_1244),
            .b(out_1512),
            .outp(out_2720)
        );        
        

        logic [WIDTH-1:0] out_2721;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2721 (
            .a(out_2720),
            .b(out_2714),
            .outp(out_2721)
        );        
        

        logic [WIDTH-1:0] out_2722;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2722 (
            .a(out_2721),
            .b(out_2717),
            .outp(out_2722)
        );        
        

        logic [WIDTH-1:0] out_2723;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2723 (
            .in(out_2714),
            .outp(out_2723)
        );
        

        logic [WIDTH-1:0] out_2724;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2724 (
            .a(out_1529),
            .b(out_2723),
            .outp(out_2724)
        );        
        

        logic [WIDTH-1:0] out_2725;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2725 (
            .in(out_2724),
            .outp(out_2725)
        );
        

        logic [WIDTH-1:0] out_2726;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2726 (
            .a(out_336),
            .b(out_2725),
            .outp(out_2726)
        );        
        

        logic [WIDTH-1:0] out_2727;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2727 (
            .a(out_2722),
            .b(out_2726),
            .outp(out_2727)
        );        
        

        logic [WIDTH-1:0] out_2728;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2728 (
            .a(out_2725),
            .b(out_343),
            .outp(out_2728)
        );        
        

        logic [WIDTH-1:0] out_2729;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2729 (
            .a(out_2727),
            .b(out_2728),
            .outp(out_2729)
        );        
        

        logic [WIDTH-1:0] out_2730;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2730 (
            .a(out_2719),
            .b(out_2729),
            .outp(out_2730)
        );        
        

        logic [WIDTH-1:0] out_2731;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2731 (
            .a(out_1244),
            .b(out_1427),
            .outp(out_2731)
        );        
        

        logic [WIDTH-1:0] out_2732;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2732 (
            .a(out_2731),
            .b(out_1355),
            .outp(out_2732)
        );        
        

        logic [WIDTH-1:0] out_2733;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.5855)
        ) inst_2733 (
            .outp(out_2733)
        );
        

        logic [WIDTH-1:0] out_2734;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2734 (
            .a(out_2733),
            .b(out_3),
            .outp(out_2734)
        );        
        

        logic [WIDTH-1:0] out_2735;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2735 (
            .a(out_2732),
            .b(out_2734),
            .outp(out_2735)
        );        
        

        logic [WIDTH-1:0] out_2736;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2736 (
            .a(out_2730),
            .b(out_2735),
            .outp(out_2736)
        );        
        

        logic [WIDTH-1:0] out_2737;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2737 (
            .a(out_1244),
            .b(out_1338),
            .outp(out_2737)
        );        
        

        logic [WIDTH-1:0] out_2738;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2355)
        ) inst_2738 (
            .outp(out_2738)
        );
        

        logic [WIDTH-1:0] out_2739;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2739 (
            .a(out_3),
            .b(out_2738),
            .outp(out_2739)
        );        
        

        logic [WIDTH-1:0] out_2740;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2740 (
            .a(out_2737),
            .b(out_2739),
            .outp(out_2740)
        );        
        

        logic [WIDTH-1:0] out_2741;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2741 (
            .a(out_2740),
            .b(out_1358),
            .outp(out_2741)
        );        
        

        logic [WIDTH-1:0] out_2742;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2742 (
            .a(out_2736),
            .b(out_2741),
            .outp(out_2742)
        );        
        

        logic [WIDTH-1:0] out_2743;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.97857)
        ) inst_2743 (
            .outp(out_2743)
        );
        

        logic [WIDTH-1:0] out_2744;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2744 (
            .a(out_2743),
            .b(out_194),
            .outp(out_2744)
        );        
        

        logic [WIDTH-1:0] out_2745;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2745 (
            .a(out_2161),
            .b(out_2744),
            .outp(out_2745)
        );        
        

        logic [WIDTH-1:0] out_2746;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(9.52857)
        ) inst_2746 (
            .outp(out_2746)
        );
        

        logic [WIDTH-1:0] out_2747;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2747 (
            .a(out_2746),
            .b(out_194),
            .outp(out_2747)
        );        
        

        logic [WIDTH-1:0] out_2748;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2748 (
            .in(out_2747),
            .outp(out_2748)
        );
        

        logic [WIDTH-1:0] out_2749;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2749 (
            .a(out_2745),
            .b(out_2748),
            .outp(out_2749)
        );        
        

        logic [WIDTH-1:0] out_2750;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(11.2232)
        ) inst_2750 (
            .outp(out_2750)
        );
        

        logic [WIDTH-1:0] out_2751;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2751 (
            .a(out_2750),
            .b(out_204),
            .outp(out_2751)
        );        
        

        logic [WIDTH-1:0] out_2752;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2752 (
            .in(out_2751),
            .outp(out_2752)
        );
        

        logic [WIDTH-1:0] out_2753;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2753 (
            .a(out_2175),
            .b(out_2752),
            .outp(out_2753)
        );        
        

        logic [WIDTH-1:0] out_2754;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2754 (
            .in(out_2753),
            .outp(out_2754)
        );
        

        logic [WIDTH-1:0] out_2755;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2755 (
            .a(out_200),
            .b(out_2754),
            .outp(out_2755)
        );        
        

        logic [WIDTH-1:0] out_2756;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2756 (
            .a(out_2749),
            .b(out_2755),
            .outp(out_2756)
        );        
        

        logic [WIDTH-1:0] out_2757;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2757 (
            .in(out_2744),
            .outp(out_2757)
        );
        

        logic [WIDTH-1:0] out_2758;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2758 (
            .a(out_2175),
            .b(out_2757),
            .outp(out_2758)
        );        
        

        logic [WIDTH-1:0] out_2759;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2759 (
            .in(out_2758),
            .outp(out_2759)
        );
        

        logic [WIDTH-1:0] out_2760;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2760 (
            .a(out_2759),
            .b(out_214),
            .outp(out_2760)
        );        
        

        logic [WIDTH-1:0] out_2761;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2761 (
            .a(out_2756),
            .b(out_2760),
            .outp(out_2761)
        );        
        

        logic [WIDTH-1:0] out_2762;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2762 (
            .a(out_2742),
            .b(out_2761),
            .outp(out_2762)
        );        
        

        logic [WIDTH-1:0] out_2763;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.79)
        ) inst_2763 (
            .outp(out_2763)
        );
        

        logic [WIDTH-1:0] out_2764;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2764 (
            .a(out_2763),
            .b(out_3),
            .outp(out_2764)
        );        
        

        logic [WIDTH-1:0] out_2765;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2765 (
            .a(out_2273),
            .b(out_2764),
            .outp(out_2765)
        );        
        

        logic [WIDTH-1:0] out_2766;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.89)
        ) inst_2766 (
            .outp(out_2766)
        );
        

        logic [WIDTH-1:0] out_2767;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2767 (
            .a(out_2766),
            .b(out_3),
            .outp(out_2767)
        );        
        

        logic [WIDTH-1:0] out_2768;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2768 (
            .in(out_2767),
            .outp(out_2768)
        );
        

        logic [WIDTH-1:0] out_2769;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2769 (
            .a(out_2765),
            .b(out_2768),
            .outp(out_2769)
        );        
        

        logic [WIDTH-1:0] out_2770;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2770 (
            .a(out_2762),
            .b(out_2769),
            .outp(out_2770)
        );        
        

        logic [WIDTH-1:0] out_2771;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.97857)
        ) inst_2771 (
            .outp(out_2771)
        );
        

        logic [WIDTH-1:0] out_2772;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2772 (
            .a(out_2771),
            .b(out_3),
            .outp(out_2772)
        );        
        

        logic [WIDTH-1:0] out_2773;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2773 (
            .a(out_2772),
            .b(out_1495),
            .outp(out_2773)
        );        
        

        logic [WIDTH-1:0] out_2774;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2774 (
            .in(out_2773),
            .outp(out_2774)
        );
        

        logic [WIDTH-1:0] out_2775;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2775 (
            .a(out_753),
            .b(out_2774),
            .outp(out_2775)
        );        
        

        logic [WIDTH-1:0] out_2776;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2776 (
            .in(out_2775),
            .outp(out_2776)
        );
        

        logic [WIDTH-1:0] out_2777;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2777 (
            .a(out_9),
            .b(out_2776),
            .outp(out_2777)
        );        
        

        logic [WIDTH-1:0] out_2778;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2778 (
            .a(out_2776),
            .b(out_21),
            .outp(out_2778)
        );        
        

        logic [WIDTH-1:0] out_2779;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2779 (
            .a(out_2777),
            .b(out_2778),
            .outp(out_2779)
        );        
        

        logic [WIDTH-1:0] out_2780;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2780 (
            .a(out_2770),
            .b(out_2779),
            .outp(out_2780)
        );        
        

        logic [WIDTH-1:0] out_2781;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.45)
        ) inst_2781 (
            .outp(out_2781)
        );
        

        logic [WIDTH-1:0] out_2782;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2782 (
            .a(out_2781),
            .b(out_3),
            .outp(out_2782)
        );        
        

        logic [WIDTH-1:0] out_2783;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2783 (
            .a(out_2315),
            .b(out_2782),
            .outp(out_2783)
        );        
        

        logic [WIDTH-1:0] out_2784;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.95)
        ) inst_2784 (
            .outp(out_2784)
        );
        

        logic [WIDTH-1:0] out_2785;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2785 (
            .a(out_2784),
            .b(out_3),
            .outp(out_2785)
        );        
        

        logic [WIDTH-1:0] out_2786;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2786 (
            .in(out_2785),
            .outp(out_2786)
        );
        

        logic [WIDTH-1:0] out_2787;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2787 (
            .a(out_2783),
            .b(out_2786),
            .outp(out_2787)
        );        
        

        logic [WIDTH-1:0] out_2788;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.725)
        ) inst_2788 (
            .outp(out_2788)
        );
        

        logic [WIDTH-1:0] out_2789;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2789 (
            .a(out_2788),
            .b(out_3),
            .outp(out_2789)
        );        
        

        logic [WIDTH-1:0] out_2790;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2790 (
            .in(out_2789),
            .outp(out_2790)
        );
        

        logic [WIDTH-1:0] out_2791;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2791 (
            .a(out_753),
            .b(out_2790),
            .outp(out_2791)
        );        
        

        logic [WIDTH-1:0] out_2792;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2792 (
            .in(out_2791),
            .outp(out_2792)
        );
        

        logic [WIDTH-1:0] out_2793;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2793 (
            .a(out_2792),
            .b(out_21),
            .outp(out_2793)
        );        
        

        logic [WIDTH-1:0] out_2794;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.42)
        ) inst_2794 (
            .outp(out_2794)
        );
        

        logic [WIDTH-1:0] out_2795;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2795 (
            .a(out_2794),
            .b(out_556),
            .outp(out_2795)
        );        
        

        logic [WIDTH-1:0] out_2796;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2796 (
            .a(out_2795),
            .b(out_559),
            .outp(out_2796)
        );        
        

        logic [WIDTH-1:0] out_2797;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2797 (
            .a(out_2290),
            .b(out_2796),
            .outp(out_2797)
        );        
        

        logic [WIDTH-1:0] out_2798;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.085)
        ) inst_2798 (
            .outp(out_2798)
        );
        

        logic [WIDTH-1:0] out_2799;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2799 (
            .a(out_2653),
            .b(out_2798),
            .outp(out_2799)
        );        
        

        logic [WIDTH-1:0] out_2800;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2800 (
            .in(out_2799),
            .outp(out_2800)
        );
        

        logic [WIDTH-1:0] out_2801;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2801 (
            .a(out_2797),
            .b(out_2800),
            .outp(out_2801)
        );        
        

        logic [WIDTH-1:0] out_2802;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.085)
        ) inst_2802 (
            .outp(out_2802)
        );
        

        logic [WIDTH-1:0] out_2803;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2803 (
            .a(out_2653),
            .b(out_2802),
            .outp(out_2803)
        );        
        

        logic [WIDTH-1:0] out_2804;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2804 (
            .a(out_2300),
            .b(out_2803),
            .outp(out_2804)
        );        
        

        logic [WIDTH-1:0] out_2805;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2805 (
            .a(out_559),
            .b(out_2795),
            .outp(out_2805)
        );        
        

        logic [WIDTH-1:0] out_2806;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2806 (
            .a(out_2804),
            .b(out_2805),
            .outp(out_2806)
        );        
        

        logic [WIDTH-1:0] out_2807;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2807 (
            .a(out_2801),
            .b(out_2806),
            .outp(out_2807)
        );        
        

        logic [WIDTH-1:0] out_2808;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2808 (
            .in(out_2807),
            .outp(out_2808)
        );
        

        logic [WIDTH-1:0] out_2809;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2809 (
            .a(out_2793),
            .b(out_2808),
            .outp(out_2809)
        );        
        

        logic [WIDTH-1:0] out_2810;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2810 (
            .a(out_9),
            .b(out_2792),
            .outp(out_2810)
        );        
        

        logic [WIDTH-1:0] out_2811;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2811 (
            .a(out_2809),
            .b(out_2810),
            .outp(out_2811)
        );        
        

        logic [WIDTH-1:0] out_2812;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2812 (
            .a(out_2787),
            .b(out_2811),
            .outp(out_2812)
        );        
        

        logic [WIDTH-1:0] out_2813;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2813 (
            .a(out_2793),
            .b(out_2812),
            .outp(out_2813)
        );        
        

        logic [WIDTH-1:0] out_2814;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2814 (
            .a(out_2780),
            .b(out_2813),
            .outp(out_2814)
        );        
        

        logic [WIDTH-1:0] out_2815;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.44223)
        ) inst_2815 (
            .outp(out_2815)
        );
        

        logic [WIDTH-1:0] out_2816;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2816 (
            .a(out_2815),
            .b(out_127),
            .outp(out_2816)
        );        
        

        logic [WIDTH-1:0] out_2817;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2817 (
            .a(out_1011),
            .b(out_2816),
            .outp(out_2817)
        );        
        

        logic [WIDTH-1:0] out_2818;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.30723)
        ) inst_2818 (
            .outp(out_2818)
        );
        

        logic [WIDTH-1:0] out_2819;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2819 (
            .a(out_2818),
            .b(out_127),
            .outp(out_2819)
        );        
        

        logic [WIDTH-1:0] out_2820;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2820 (
            .a(out_2819),
            .b(out_1017),
            .outp(out_2820)
        );        
        

        logic [WIDTH-1:0] out_2821;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2821 (
            .a(out_2817),
            .b(out_2820),
            .outp(out_2821)
        );        
        

        logic [WIDTH-1:0] out_2822;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.08)
        ) inst_2822 (
            .outp(out_2822)
        );
        

        logic [WIDTH-1:0] out_2823;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2823 (
            .a(out_2822),
            .b(out_137),
            .outp(out_2823)
        );        
        

        logic [WIDTH-1:0] out_2824;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2824 (
            .a(out_2821),
            .b(out_2823),
            .outp(out_2824)
        );        
        

        logic [WIDTH-1:0] out_2825;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2825 (
            .a(out_2814),
            .b(out_2824),
            .outp(out_2825)
        );        
        

        logic [WIDTH-1:0] out_2826;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2826 (
            .a(out_2816),
            .b(out_1011),
            .outp(out_2826)
        );        
        

        logic [WIDTH-1:0] out_2827;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2827 (
            .in(out_2823),
            .outp(out_2827)
        );
        

        logic [WIDTH-1:0] out_2828;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2828 (
            .a(out_2826),
            .b(out_2827),
            .outp(out_2828)
        );        
        

        logic [WIDTH-1:0] out_2829;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2829 (
            .a(out_1017),
            .b(out_2819),
            .outp(out_2829)
        );        
        

        logic [WIDTH-1:0] out_2830;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2830 (
            .a(out_2828),
            .b(out_2829),
            .outp(out_2830)
        );        
        

        logic [WIDTH-1:0] out_2831;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2831 (
            .a(out_2825),
            .b(out_2830),
            .outp(out_2831)
        );        
        

        logic [WIDTH-1:0] out_2832;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2832 (
            .a(out_2822),
            .b(out_152),
            .outp(out_2832)
        );        
        

        logic [WIDTH-1:0] out_2833;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2833 (
            .in(out_2832),
            .outp(out_2833)
        );
        

        logic [WIDTH-1:0] out_2834;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.36223)
        ) inst_2834 (
            .outp(out_2834)
        );
        

        logic [WIDTH-1:0] out_2835;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2835 (
            .a(out_2834),
            .b(out_127),
            .outp(out_2835)
        );        
        

        logic [WIDTH-1:0] out_2836;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2836 (
            .a(out_1017),
            .b(out_2835),
            .outp(out_2836)
        );        
        

        logic [WIDTH-1:0] out_2837;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2837 (
            .a(out_2833),
            .b(out_2836),
            .outp(out_2837)
        );        
        

        logic [WIDTH-1:0] out_2838;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.38723)
        ) inst_2838 (
            .outp(out_2838)
        );
        

        logic [WIDTH-1:0] out_2839;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2839 (
            .a(out_2838),
            .b(out_127),
            .outp(out_2839)
        );        
        

        logic [WIDTH-1:0] out_2840;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2840 (
            .a(out_2839),
            .b(out_1011),
            .outp(out_2840)
        );        
        

        logic [WIDTH-1:0] out_2841;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2841 (
            .a(out_2837),
            .b(out_2840),
            .outp(out_2841)
        );        
        

        logic [WIDTH-1:0] out_2842;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2842 (
            .a(out_2831),
            .b(out_2841),
            .outp(out_2842)
        );        
        

        logic [WIDTH-1:0] out_2843;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2843 (
            .a(out_2835),
            .b(out_1017),
            .outp(out_2843)
        );        
        

        logic [WIDTH-1:0] out_2844;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2844 (
            .a(out_2832),
            .b(out_2843),
            .outp(out_2844)
        );        
        

        logic [WIDTH-1:0] out_2845;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2845 (
            .a(out_1011),
            .b(out_2839),
            .outp(out_2845)
        );        
        

        logic [WIDTH-1:0] out_2846;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2846 (
            .a(out_2844),
            .b(out_2845),
            .outp(out_2846)
        );        
        

        logic [WIDTH-1:0] out_2847;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2847 (
            .a(out_2842),
            .b(out_2846),
            .outp(out_2847)
        );        
        

        logic [WIDTH-1:0] out_2848;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2848 (
            .a(out_2817),
            .b(out_2843),
            .outp(out_2848)
        );        
        

        logic [WIDTH-1:0] out_2849;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.025)
        ) inst_2849 (
            .outp(out_2849)
        );
        

        logic [WIDTH-1:0] out_2850;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2850 (
            .a(out_2849),
            .b(out_137),
            .outp(out_2850)
        );        
        

        logic [WIDTH-1:0] out_2851;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2851 (
            .a(out_2848),
            .b(out_2850),
            .outp(out_2851)
        );        
        

        logic [WIDTH-1:0] out_2852;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2852 (
            .a(out_2847),
            .b(out_2851),
            .outp(out_2852)
        );        
        

        logic [WIDTH-1:0] out_2853;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2853 (
            .a(out_2826),
            .b(out_2836),
            .outp(out_2853)
        );        
        

        logic [WIDTH-1:0] out_2854;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2854 (
            .in(out_2850),
            .outp(out_2854)
        );
        

        logic [WIDTH-1:0] out_2855;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2855 (
            .a(out_2853),
            .b(out_2854),
            .outp(out_2855)
        );        
        

        logic [WIDTH-1:0] out_2856;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2856 (
            .a(out_2852),
            .b(out_2855),
            .outp(out_2856)
        );        
        

        logic [WIDTH-1:0] out_2857;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.80223)
        ) inst_2857 (
            .outp(out_2857)
        );
        

        logic [WIDTH-1:0] out_2858;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2858 (
            .a(out_2857),
            .b(out_1011),
            .outp(out_2858)
        );        
        

        logic [WIDTH-1:0] out_2859;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2859 (
            .a(out_2858),
            .b(out_127),
            .outp(out_2859)
        );        
        

        logic [WIDTH-1:0] out_2860;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2860 (
            .in(out_2859),
            .outp(out_2860)
        );
        

        logic [WIDTH-1:0] out_2861;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2861 (
            .a(out_2833),
            .b(out_2860),
            .outp(out_2861)
        );        
        

        logic [WIDTH-1:0] out_2862;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.82723)
        ) inst_2862 (
            .outp(out_2862)
        );
        

        logic [WIDTH-1:0] out_2863;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2863 (
            .a(out_2862),
            .b(out_1017),
            .outp(out_2863)
        );        
        

        logic [WIDTH-1:0] out_2864;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2864 (
            .a(out_2863),
            .b(out_127),
            .outp(out_2864)
        );        
        

        logic [WIDTH-1:0] out_2865;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2865 (
            .a(out_2861),
            .b(out_2864),
            .outp(out_2865)
        );        
        

        logic [WIDTH-1:0] out_2866;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2866 (
            .a(out_2856),
            .b(out_2865),
            .outp(out_2866)
        );        
        

        logic [WIDTH-1:0] out_2867;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2867 (
            .a(out_2832),
            .b(out_2859),
            .outp(out_2867)
        );        
        

        logic [WIDTH-1:0] out_2868;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2868 (
            .in(out_2864),
            .outp(out_2868)
        );
        

        logic [WIDTH-1:0] out_2869;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2869 (
            .a(out_2867),
            .b(out_2868),
            .outp(out_2869)
        );        
        

        logic [WIDTH-1:0] out_2870;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2870 (
            .a(out_2866),
            .b(out_2869),
            .outp(out_2870)
        );        
        

        logic [WIDTH-1:0] out_2871;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2871 (
            .a(out_2850),
            .b(out_2868),
            .outp(out_2871)
        );        
        

        logic [WIDTH-1:0] out_2872;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.74723)
        ) inst_2872 (
            .outp(out_2872)
        );
        

        logic [WIDTH-1:0] out_2873;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2873 (
            .a(out_2872),
            .b(out_1011),
            .outp(out_2873)
        );        
        

        logic [WIDTH-1:0] out_2874;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2874 (
            .a(out_2873),
            .b(out_127),
            .outp(out_2874)
        );        
        

        logic [WIDTH-1:0] out_2875;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2875 (
            .a(out_2871),
            .b(out_2874),
            .outp(out_2875)
        );        
        

        logic [WIDTH-1:0] out_2876;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2876 (
            .a(out_2870),
            .b(out_2875),
            .outp(out_2876)
        );        
        

        logic [WIDTH-1:0] out_2877;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2877 (
            .a(out_2854),
            .b(out_2864),
            .outp(out_2877)
        );        
        

        logic [WIDTH-1:0] out_2878;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2878 (
            .in(out_2874),
            .outp(out_2878)
        );
        

        logic [WIDTH-1:0] out_2879;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2879 (
            .a(out_2877),
            .b(out_2878),
            .outp(out_2879)
        );        
        

        logic [WIDTH-1:0] out_2880;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2880 (
            .a(out_2876),
            .b(out_2879),
            .outp(out_2880)
        );        
        

        logic [WIDTH-1:0] out_2881;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.5325)
        ) inst_2881 (
            .outp(out_2881)
        );
        

        logic [WIDTH-1:0] out_2882;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2882 (
            .a(out_2881),
            .b(out_3),
            .outp(out_2882)
        );        
        

        logic [WIDTH-1:0] out_2883;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6325)
        ) inst_2883 (
            .outp(out_2883)
        );
        

        logic [WIDTH-1:0] out_2884;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2884 (
            .a(out_2883),
            .b(out_3),
            .outp(out_2884)
        );        
        

        logic [WIDTH-1:0] out_2885;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2885 (
            .in(out_2884),
            .outp(out_2885)
        );
        

        logic [WIDTH-1:0] out_2886;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2886 (
            .a(out_2882),
            .b(out_2885),
            .outp(out_2886)
        );        
        

        logic [WIDTH-1:0] out_2887;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.25)
        ) inst_2887 (
            .outp(out_2887)
        );
        

        logic [WIDTH-1:0] out_2888;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2888 (
            .a(out_2887),
            .b(out_14),
            .outp(out_2888)
        );        
        

        logic [WIDTH-1:0] out_2889;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2889 (
            .a(out_2886),
            .b(out_2888),
            .outp(out_2889)
        );        
        

        logic [WIDTH-1:0] out_2890;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.8)
        ) inst_2890 (
            .outp(out_2890)
        );
        

        logic [WIDTH-1:0] out_2891;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2891 (
            .a(out_2890),
            .b(out_14),
            .outp(out_2891)
        );        
        

        logic [WIDTH-1:0] out_2892;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2892 (
            .in(out_2891),
            .outp(out_2892)
        );
        

        logic [WIDTH-1:0] out_2893;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2893 (
            .a(out_2889),
            .b(out_2892),
            .outp(out_2893)
        );        
        

        logic [WIDTH-1:0] out_2894;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2894 (
            .a(out_2880),
            .b(out_2893),
            .outp(out_2894)
        );        
        

        logic [WIDTH-1:0] out_2895;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.63929)
        ) inst_2895 (
            .outp(out_2895)
        );
        

        logic [WIDTH-1:0] out_2896;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2896 (
            .a(out_2895),
            .b(out_194),
            .outp(out_2896)
        );        
        

        logic [WIDTH-1:0] out_2897;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.18929)
        ) inst_2897 (
            .outp(out_2897)
        );
        

        logic [WIDTH-1:0] out_2898;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2898 (
            .a(out_2897),
            .b(out_194),
            .outp(out_2898)
        );        
        

        logic [WIDTH-1:0] out_2899;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2899 (
            .in(out_2898),
            .outp(out_2899)
        );
        

        logic [WIDTH-1:0] out_2900;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2900 (
            .a(out_2896),
            .b(out_2899),
            .outp(out_2900)
        );        
        

        logic [WIDTH-1:0] out_2901;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.79911)
        ) inst_2901 (
            .outp(out_2901)
        );
        

        logic [WIDTH-1:0] out_2902;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2902 (
            .a(out_2901),
            .b(out_204),
            .outp(out_2902)
        );        
        

        logic [WIDTH-1:0] out_2903;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2903 (
            .in(out_2902),
            .outp(out_2903)
        );
        

        logic [WIDTH-1:0] out_2904;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2904 (
            .in(out_2891),
            .outp(out_2904)
        );
        

        logic [WIDTH-1:0] out_2905;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2905 (
            .a(out_2903),
            .b(out_2904),
            .outp(out_2905)
        );        
        

        logic [WIDTH-1:0] out_2906;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2906 (
            .in(out_2905),
            .outp(out_2906)
        );
        

        logic [WIDTH-1:0] out_2907;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2907 (
            .a(out_200),
            .b(out_2906),
            .outp(out_2907)
        );        
        

        logic [WIDTH-1:0] out_2908;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2908 (
            .a(out_2900),
            .b(out_2907),
            .outp(out_2908)
        );        
        

        logic [WIDTH-1:0] out_2909;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2909 (
            .in(out_2896),
            .outp(out_2909)
        );
        

        logic [WIDTH-1:0] out_2910;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2910 (
            .a(out_2909),
            .b(out_2904),
            .outp(out_2910)
        );        
        

        logic [WIDTH-1:0] out_2911;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2911 (
            .in(out_2910),
            .outp(out_2911)
        );
        

        logic [WIDTH-1:0] out_2912;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2912 (
            .a(out_2911),
            .b(out_214),
            .outp(out_2912)
        );        
        

        logic [WIDTH-1:0] out_2913;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2913 (
            .a(out_2908),
            .b(out_2912),
            .outp(out_2913)
        );        
        

        logic [WIDTH-1:0] out_2914;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2914 (
            .a(out_2913),
            .b(out_2888),
            .outp(out_2914)
        );        
        

        logic [WIDTH-1:0] out_2915;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2915 (
            .a(out_2914),
            .b(out_2892),
            .outp(out_2915)
        );        
        

        logic [WIDTH-1:0] out_2916;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2916 (
            .a(out_2894),
            .b(out_2915),
            .outp(out_2916)
        );        
        

        logic [WIDTH-1:0] out_2917;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.7575)
        ) inst_2917 (
            .outp(out_2917)
        );
        

        logic [WIDTH-1:0] out_2918;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2918 (
            .a(out_2917),
            .b(out_3),
            .outp(out_2918)
        );        
        

        logic [WIDTH-1:0] out_2919;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.8575)
        ) inst_2919 (
            .outp(out_2919)
        );
        

        logic [WIDTH-1:0] out_2920;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2920 (
            .a(out_2919),
            .b(out_3),
            .outp(out_2920)
        );        
        

        logic [WIDTH-1:0] out_2921;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2921 (
            .in(out_2920),
            .outp(out_2921)
        );
        

        logic [WIDTH-1:0] out_2922;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2922 (
            .a(out_2918),
            .b(out_2921),
            .outp(out_2922)
        );        
        

        logic [WIDTH-1:0] out_2923;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2923 (
            .a(out_2922),
            .b(out_2888),
            .outp(out_2923)
        );        
        

        logic [WIDTH-1:0] out_2924;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2924 (
            .a(out_2923),
            .b(out_2892),
            .outp(out_2924)
        );        
        

        logic [WIDTH-1:0] out_2925;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2925 (
            .a(out_2916),
            .b(out_2924),
            .outp(out_2925)
        );        
        

        logic [WIDTH-1:0] out_2926;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.8075)
        ) inst_2926 (
            .outp(out_2926)
        );
        

        logic [WIDTH-1:0] out_2927;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2927 (
            .a(out_2926),
            .b(out_3),
            .outp(out_2927)
        );        
        

        logic [WIDTH-1:0] out_2928;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2928 (
            .in(out_2927),
            .outp(out_2928)
        );
        

        logic [WIDTH-1:0] out_2929;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0999999)
        ) inst_2929 (
            .outp(out_2929)
        );
        

        logic [WIDTH-1:0] out_2930;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2930 (
            .a(out_2929),
            .b(out_14),
            .outp(out_2930)
        );        
        

        logic [WIDTH-1:0] out_2931;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2931 (
            .in(out_2930),
            .outp(out_2931)
        );
        

        logic [WIDTH-1:0] out_2932;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2932 (
            .a(out_2928),
            .b(out_2931),
            .outp(out_2932)
        );        
        

        logic [WIDTH-1:0] out_2933;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2933 (
            .in(out_2932),
            .outp(out_2933)
        );
        

        logic [WIDTH-1:0] out_2934;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2934 (
            .a(out_2933),
            .b(out_460),
            .outp(out_2934)
        );        
        

        logic [WIDTH-1:0] out_2935;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2935 (
            .a(out_2925),
            .b(out_2934),
            .outp(out_2935)
        );        
        

        logic [WIDTH-1:0] out_2936;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.0025)
        ) inst_2936 (
            .outp(out_2936)
        );
        

        logic [WIDTH-1:0] out_2937;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2937 (
            .a(out_2936),
            .b(out_3),
            .outp(out_2937)
        );        
        

        logic [WIDTH-1:0] out_2938;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.1025)
        ) inst_2938 (
            .outp(out_2938)
        );
        

        logic [WIDTH-1:0] out_2939;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2939 (
            .a(out_2938),
            .b(out_3),
            .outp(out_2939)
        );        
        

        logic [WIDTH-1:0] out_2940;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2940 (
            .in(out_2939),
            .outp(out_2940)
        );
        

        logic [WIDTH-1:0] out_2941;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2941 (
            .a(out_2937),
            .b(out_2940),
            .outp(out_2941)
        );        
        

        logic [WIDTH-1:0] out_2942;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2942 (
            .a(out_2941),
            .b(out_2892),
            .outp(out_2942)
        );        
        

        logic [WIDTH-1:0] out_2943;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.45)
        ) inst_2943 (
            .outp(out_2943)
        );
        

        logic [WIDTH-1:0] out_2944;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2944 (
            .a(out_2943),
            .b(out_14),
            .outp(out_2944)
        );        
        

        logic [WIDTH-1:0] out_2945;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2945 (
            .a(out_2942),
            .b(out_2944),
            .outp(out_2945)
        );        
        

        logic [WIDTH-1:0] out_2946;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2946 (
            .a(out_2935),
            .b(out_2945),
            .outp(out_2946)
        );        
        

        logic [WIDTH-1:0] out_2947;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0154991)
        ) inst_2947 (
            .outp(out_2947)
        );
        

        logic [WIDTH-1:0] out_2948;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2948 (
            .a(out_3),
            .b(out_2947),
            .outp(out_2948)
        );        
        

        logic [WIDTH-1:0] out_2949;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.084501)
        ) inst_2949 (
            .outp(out_2949)
        );
        

        logic [WIDTH-1:0] out_2950;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2950 (
            .a(out_2949),
            .b(out_3),
            .outp(out_2950)
        );        
        

        logic [WIDTH-1:0] out_2951;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2951 (
            .in(out_2950),
            .outp(out_2951)
        );
        

        logic [WIDTH-1:0] out_2952;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2952 (
            .a(out_2948),
            .b(out_2951),
            .outp(out_2952)
        );        
        

        logic [WIDTH-1:0] out_2953;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2953 (
            .a(out_2952),
            .b(out_2892),
            .outp(out_2953)
        );        
        

        logic [WIDTH-1:0] out_2954;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2954 (
            .a(out_2953),
            .b(out_2944),
            .outp(out_2954)
        );        
        

        logic [WIDTH-1:0] out_2955;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2955 (
            .a(out_2946),
            .b(out_2954),
            .outp(out_2955)
        );        
        

        logic [WIDTH-1:0] out_2956;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.11593)
        ) inst_2956 (
            .outp(out_2956)
        );
        

        logic [WIDTH-1:0] out_2957;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2957 (
            .a(out_2956),
            .b(out_3),
            .outp(out_2957)
        );        
        

        logic [WIDTH-1:0] out_2958;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2958 (
            .a(out_2957),
            .b(out_1495),
            .outp(out_2958)
        );        
        

        logic [WIDTH-1:0] out_2959;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2959 (
            .in(out_2958),
            .outp(out_2959)
        );
        

        logic [WIDTH-1:0] out_2960;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.525)
        ) inst_2960 (
            .outp(out_2960)
        );
        

        logic [WIDTH-1:0] out_2961;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2961 (
            .a(out_2960),
            .b(out_14),
            .outp(out_2961)
        );        
        

        logic [WIDTH-1:0] out_2962;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2962 (
            .in(out_2961),
            .outp(out_2962)
        );
        

        logic [WIDTH-1:0] out_2963;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2963 (
            .a(out_2959),
            .b(out_2962),
            .outp(out_2963)
        );        
        

        logic [WIDTH-1:0] out_2964;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2964 (
            .in(out_2963),
            .outp(out_2964)
        );
        

        logic [WIDTH-1:0] out_2965;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2965 (
            .a(out_9),
            .b(out_2964),
            .outp(out_2965)
        );        
        

        logic [WIDTH-1:0] out_2966;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2966 (
            .a(out_2964),
            .b(out_21),
            .outp(out_2966)
        );        
        

        logic [WIDTH-1:0] out_2967;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2967 (
            .a(out_2965),
            .b(out_2966),
            .outp(out_2967)
        );        
        

        logic [WIDTH-1:0] out_2968;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2968 (
            .a(out_2955),
            .b(out_2967),
            .outp(out_2968)
        );        
        

        logic [WIDTH-1:0] out_2969;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6945)
        ) inst_2969 (
            .outp(out_2969)
        );
        

        logic [WIDTH-1:0] out_2970;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2970 (
            .a(out_2969),
            .b(out_3),
            .outp(out_2970)
        );        
        

        logic [WIDTH-1:0] out_2971;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.794501)
        ) inst_2971 (
            .outp(out_2971)
        );
        

        logic [WIDTH-1:0] out_2972;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2972 (
            .a(out_2971),
            .b(out_3),
            .outp(out_2972)
        );        
        

        logic [WIDTH-1:0] out_2973;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2973 (
            .in(out_2972),
            .outp(out_2973)
        );
        

        logic [WIDTH-1:0] out_2974;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2974 (
            .a(out_2970),
            .b(out_2973),
            .outp(out_2974)
        );        
        

        logic [WIDTH-1:0] out_2975;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2975 (
            .a(out_2974),
            .b(out_2961),
            .outp(out_2975)
        );        
        

        logic [WIDTH-1:0] out_2976;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2976 (
            .a(out_2975),
            .b(out_2892),
            .outp(out_2976)
        );        
        

        logic [WIDTH-1:0] out_2977;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2977 (
            .a(out_2968),
            .b(out_2976),
            .outp(out_2977)
        );        
        

        logic [WIDTH-1:0] out_2978;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.1445)
        ) inst_2978 (
            .outp(out_2978)
        );
        

        logic [WIDTH-1:0] out_2979;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2979 (
            .a(out_2978),
            .b(out_3),
            .outp(out_2979)
        );        
        

        logic [WIDTH-1:0] out_2980;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2445)
        ) inst_2980 (
            .outp(out_2980)
        );
        

        logic [WIDTH-1:0] out_2981;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2981 (
            .a(out_2980),
            .b(out_3),
            .outp(out_2981)
        );        
        

        logic [WIDTH-1:0] out_2982;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2982 (
            .in(out_2981),
            .outp(out_2982)
        );
        

        logic [WIDTH-1:0] out_2983;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2983 (
            .a(out_2979),
            .b(out_2982),
            .outp(out_2983)
        );        
        

        logic [WIDTH-1:0] out_2984;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.2)
        ) inst_2984 (
            .outp(out_2984)
        );
        

        logic [WIDTH-1:0] out_2985;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2985 (
            .a(out_14),
            .b(out_2984),
            .outp(out_2985)
        );        
        

        logic [WIDTH-1:0] out_2986;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2986 (
            .a(out_2983),
            .b(out_2985),
            .outp(out_2986)
        );        
        

        logic [WIDTH-1:0] out_2987;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2987 (
            .a(out_2986),
            .b(out_2892),
            .outp(out_2987)
        );        
        

        logic [WIDTH-1:0] out_2988;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2988 (
            .a(out_2977),
            .b(out_2987),
            .outp(out_2988)
        );        
        

        logic [WIDTH-1:0] out_2989;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2989 (
            .a(out_2970),
            .b(out_2982),
            .outp(out_2989)
        );        
        

        logic [WIDTH-1:0] out_2990;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.525)
        ) inst_2990 (
            .outp(out_2990)
        );
        

        logic [WIDTH-1:0] out_2991;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2991 (
            .a(out_2990),
            .b(out_14),
            .outp(out_2991)
        );        
        

        logic [WIDTH-1:0] out_2992;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2992 (
            .in(out_2991),
            .outp(out_2992)
        );
        

        logic [WIDTH-1:0] out_2993;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2993 (
            .a(out_2989),
            .b(out_2992),
            .outp(out_2993)
        );        
        

        logic [WIDTH-1:0] out_2994;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.969501)
        ) inst_2994 (
            .outp(out_2994)
        );
        

        logic [WIDTH-1:0] out_2995;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2995 (
            .a(out_2994),
            .b(out_3),
            .outp(out_2995)
        );        
        

        logic [WIDTH-1:0] out_2996;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2996 (
            .in(out_2995),
            .outp(out_2996)
        );
        

        logic [WIDTH-1:0] out_2997;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2997 (
            .a(out_2996),
            .b(out_2962),
            .outp(out_2997)
        );        
        

        logic [WIDTH-1:0] out_2998;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2998 (
            .in(out_2997),
            .outp(out_2998)
        );
        

        logic [WIDTH-1:0] out_2999;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_2999 (
            .a(out_9),
            .b(out_2998),
            .outp(out_2999)
        );        
        

        logic [WIDTH-1:0] out_3000;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3000 (
            .a(out_2993),
            .b(out_2999),
            .outp(out_3000)
        );        
        

        logic [WIDTH-1:0] out_3001;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3001 (
            .a(out_2998),
            .b(out_21),
            .outp(out_3001)
        );        
        

        logic [WIDTH-1:0] out_3002;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3002 (
            .a(out_3000),
            .b(out_3001),
            .outp(out_3002)
        );        
        

        logic [WIDTH-1:0] out_3003;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3003 (
            .a(out_3002),
            .b(out_2888),
            .outp(out_3003)
        );        
        

        logic [WIDTH-1:0] out_3004;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3004 (
            .a(out_2988),
            .b(out_3003),
            .outp(out_3004)
        );        
        

        logic [WIDTH-1:0] out_3005;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.289485)
        ) inst_3005 (
            .outp(out_3005)
        );
        

        logic [WIDTH-1:0] out_3006;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3006 (
            .a(out_3005),
            .b(out_1826),
            .outp(out_3006)
        );        
        

        logic [WIDTH-1:0] out_3007;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3007 (
            .a(out_1823),
            .b(out_3006),
            .outp(out_3007)
        );        
        

        logic [WIDTH-1:0] out_3008;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.707348)
        ) inst_3008 (
            .outp(out_3008)
        );
        

        logic [WIDTH-1:0] out_3009;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3009 (
            .a(out_3008),
            .b(out_1831),
            .outp(out_3009)
        );        
        

        logic [WIDTH-1:0] out_3010;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3010 (
            .a(out_3007),
            .b(out_3009),
            .outp(out_3010)
        );        
        

        logic [WIDTH-1:0] out_3011;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.570488)
        ) inst_3011 (
            .outp(out_3011)
        );
        

        logic [WIDTH-1:0] out_3012;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3012 (
            .a(out_3011),
            .b(out_1834),
            .outp(out_3012)
        );        
        

        logic [WIDTH-1:0] out_3013;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3013 (
            .in(out_3012),
            .outp(out_3013)
        );
        

        logic [WIDTH-1:0] out_3014;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3014 (
            .a(out_3010),
            .b(out_3013),
            .outp(out_3014)
        );        
        

        logic [WIDTH-1:0] out_3015;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3015 (
            .in(out_3009),
            .outp(out_3015)
        );
        

        logic [WIDTH-1:0] out_3016;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3016 (
            .a(out_3012),
            .b(out_3015),
            .outp(out_3016)
        );        
        

        logic [WIDTH-1:0] out_3017;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3017 (
            .a(out_3006),
            .b(out_1823),
            .outp(out_3017)
        );        
        

        logic [WIDTH-1:0] out_3018;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3018 (
            .a(out_3016),
            .b(out_3017),
            .outp(out_3018)
        );        
        

        logic [WIDTH-1:0] out_3019;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3019 (
            .a(out_3014),
            .b(out_3018),
            .outp(out_3019)
        );        
        

        logic [WIDTH-1:0] out_3020;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3020 (
            .in(out_3019),
            .outp(out_3020)
        );
        

        logic [WIDTH-1:0] out_3021;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5495)
        ) inst_3021 (
            .outp(out_3021)
        );
        

        logic [WIDTH-1:0] out_3022;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3022 (
            .a(out_3021),
            .b(out_3),
            .outp(out_3022)
        );        
        

        logic [WIDTH-1:0] out_3023;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3023 (
            .in(out_3022),
            .outp(out_3023)
        );
        

        logic [WIDTH-1:0] out_3024;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3024 (
            .a(out_3023),
            .b(out_2962),
            .outp(out_3024)
        );        
        

        logic [WIDTH-1:0] out_3025;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3025 (
            .in(out_3024),
            .outp(out_3025)
        );
        

        logic [WIDTH-1:0] out_3026;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3026 (
            .a(out_9),
            .b(out_3025),
            .outp(out_3026)
        );        
        

        logic [WIDTH-1:0] out_3027;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3027 (
            .a(out_3020),
            .b(out_3026),
            .outp(out_3027)
        );        
        

        logic [WIDTH-1:0] out_3028;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3028 (
            .a(out_3025),
            .b(out_21),
            .outp(out_3028)
        );        
        

        logic [WIDTH-1:0] out_3029;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3029 (
            .a(out_3027),
            .b(out_3028),
            .outp(out_3029)
        );        
        

        logic [WIDTH-1:0] out_3030;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3030 (
            .a(out_3004),
            .b(out_3029),
            .outp(out_3030)
        );        
        

        logic [WIDTH-1:0] out_3031;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.135)
        ) inst_3031 (
            .outp(out_3031)
        );
        

        logic [WIDTH-1:0] out_3032;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3032 (
            .a(out_3031),
            .b(out_152),
            .outp(out_3032)
        );        
        

        logic [WIDTH-1:0] out_3033;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3033 (
            .in(out_3032),
            .outp(out_3033)
        );
        

        logic [WIDTH-1:0] out_3034;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3034 (
            .a(out_3033),
            .b(out_2840),
            .outp(out_3034)
        );        
        

        logic [WIDTH-1:0] out_3035;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3035 (
            .a(out_3034),
            .b(out_2829),
            .outp(out_3035)
        );        
        

        logic [WIDTH-1:0] out_3036;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3036 (
            .a(out_3030),
            .b(out_3035),
            .outp(out_3036)
        );        
        

        logic [WIDTH-1:0] out_3037;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3037 (
            .a(out_3032),
            .b(out_2820),
            .outp(out_3037)
        );        
        

        logic [WIDTH-1:0] out_3038;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3038 (
            .a(out_3037),
            .b(out_2845),
            .outp(out_3038)
        );        
        

        logic [WIDTH-1:0] out_3039;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3039 (
            .a(out_3036),
            .b(out_3038),
            .outp(out_3039)
        );        
        

        logic [WIDTH-1:0] out_3040;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.25)
        ) inst_3040 (
            .outp(out_3040)
        );
        

        logic [WIDTH-1:0] out_3041;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3041 (
            .a(out_3040),
            .b(out_3),
            .outp(out_3041)
        );        
        

        logic [WIDTH-1:0] out_3042;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3042 (
            .a(out_2992),
            .b(out_3041),
            .outp(out_3042)
        );        
        

        logic [WIDTH-1:0] out_3043;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.8)
        ) inst_3043 (
            .outp(out_3043)
        );
        

        logic [WIDTH-1:0] out_3044;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3044 (
            .a(out_3043),
            .b(out_3),
            .outp(out_3044)
        );        
        

        logic [WIDTH-1:0] out_3045;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3045 (
            .in(out_3044),
            .outp(out_3045)
        );
        

        logic [WIDTH-1:0] out_3046;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3046 (
            .a(out_3042),
            .b(out_3045),
            .outp(out_3046)
        );        
        

        logic [WIDTH-1:0] out_3047;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.525)
        ) inst_3047 (
            .outp(out_3047)
        );
        

        logic [WIDTH-1:0] out_3048;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3048 (
            .a(out_3047),
            .b(out_3),
            .outp(out_3048)
        );        
        

        logic [WIDTH-1:0] out_3049;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3049 (
            .in(out_3048),
            .outp(out_3049)
        );
        

        logic [WIDTH-1:0] out_3050;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3050 (
            .a(out_3049),
            .b(out_2962),
            .outp(out_3050)
        );        
        

        logic [WIDTH-1:0] out_3051;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3051 (
            .in(out_3050),
            .outp(out_3051)
        );
        

        logic [WIDTH-1:0] out_3052;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3052 (
            .a(out_9),
            .b(out_3051),
            .outp(out_3052)
        );        
        

        logic [WIDTH-1:0] out_3053;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3053 (
            .a(out_3046),
            .b(out_3052),
            .outp(out_3053)
        );        
        

        logic [WIDTH-1:0] out_3054;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3054 (
            .a(out_3051),
            .b(out_21),
            .outp(out_3054)
        );        
        

        logic [WIDTH-1:0] out_3055;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3055 (
            .a(out_3053),
            .b(out_3054),
            .outp(out_3055)
        );        
        

        logic [WIDTH-1:0] out_3056;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3056 (
            .a(out_3055),
            .b(out_2888),
            .outp(out_3056)
        );        
        

        logic [WIDTH-1:0] out_3057;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3057 (
            .a(out_3039),
            .b(out_3056),
            .outp(out_3057)
        );        
        

        logic [WIDTH-1:0] out_3058;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.55)
        ) inst_3058 (
            .outp(out_3058)
        );
        

        logic [WIDTH-1:0] out_3059;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3059 (
            .a(out_3058),
            .b(out_14),
            .outp(out_3059)
        );        
        

        logic [WIDTH-1:0] out_3060;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3060 (
            .in(out_3059),
            .outp(out_3060)
        );
        

        logic [WIDTH-1:0] out_3061;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.05)
        ) inst_3061 (
            .outp(out_3061)
        );
        

        logic [WIDTH-1:0] out_3062;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3062 (
            .a(out_3061),
            .b(out_3),
            .outp(out_3062)
        );        
        

        logic [WIDTH-1:0] out_3063;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3063 (
            .a(out_3060),
            .b(out_3062),
            .outp(out_3063)
        );        
        

        logic [WIDTH-1:0] out_3064;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.15)
        ) inst_3064 (
            .outp(out_3064)
        );
        

        logic [WIDTH-1:0] out_3065;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3065 (
            .a(out_3064),
            .b(out_3),
            .outp(out_3065)
        );        
        

        logic [WIDTH-1:0] out_3066;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3066 (
            .in(out_3065),
            .outp(out_3066)
        );
        

        logic [WIDTH-1:0] out_3067;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3067 (
            .a(out_3063),
            .b(out_3066),
            .outp(out_3067)
        );        
        

        logic [WIDTH-1:0] out_3068;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3068 (
            .a(out_3067),
            .b(out_2985),
            .outp(out_3068)
        );        
        

        logic [WIDTH-1:0] out_3069;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3069 (
            .a(out_3057),
            .b(out_3068),
            .outp(out_3069)
        );        
        

        logic [WIDTH-1:0] out_3070;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.9)
        ) inst_3070 (
            .outp(out_3070)
        );
        

        logic [WIDTH-1:0] out_3071;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3071 (
            .a(out_3070),
            .b(out_3),
            .outp(out_3071)
        );        
        

        logic [WIDTH-1:0] out_3072;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.3)
        ) inst_3072 (
            .outp(out_3072)
        );
        

        logic [WIDTH-1:0] out_3073;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3073 (
            .a(out_3072),
            .b(out_3),
            .outp(out_3073)
        );        
        

        logic [WIDTH-1:0] out_3074;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3074 (
            .in(out_3073),
            .outp(out_3074)
        );
        

        logic [WIDTH-1:0] out_3075;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3075 (
            .a(out_3071),
            .b(out_3074),
            .outp(out_3075)
        );        
        

        logic [WIDTH-1:0] out_3076;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.25)
        ) inst_3076 (
            .outp(out_3076)
        );
        

        logic [WIDTH-1:0] out_3077;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3077 (
            .a(out_3076),
            .b(out_14),
            .outp(out_3077)
        );        
        

        logic [WIDTH-1:0] out_3078;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3078 (
            .in(out_3077),
            .outp(out_3078)
        );
        

        logic [WIDTH-1:0] out_3079;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3079 (
            .a(out_3075),
            .b(out_3078),
            .outp(out_3079)
        );        
        

        logic [WIDTH-1:0] out_3080;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.15)
        ) inst_3080 (
            .outp(out_3080)
        );
        

        logic [WIDTH-1:0] out_3081;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3081 (
            .a(out_3080),
            .b(out_14),
            .outp(out_3081)
        );        
        

        logic [WIDTH-1:0] out_3082;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3082 (
            .a(out_3079),
            .b(out_3081),
            .outp(out_3082)
        );        
        

        logic [WIDTH-1:0] out_3083;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3083 (
            .a(out_3069),
            .b(out_3082),
            .outp(out_3083)
        );        
        

        logic [WIDTH-1:0] out_3084;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3084 (
            .a(out_3059),
            .b(out_3071),
            .outp(out_3084)
        );        
        

        logic [WIDTH-1:0] out_3085;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3085 (
            .a(out_3084),
            .b(out_3074),
            .outp(out_3085)
        );        
        

        logic [WIDTH-1:0] out_3086;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3086 (
            .in(out_3059),
            .outp(out_3086)
        );
        

        logic [WIDTH-1:0] out_3087;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3087 (
            .in(out_3071),
            .outp(out_3087)
        );
        

        logic [WIDTH-1:0] out_3088;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3088 (
            .a(out_3086),
            .b(out_3087),
            .outp(out_3088)
        );        
        

        logic [WIDTH-1:0] out_3089;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3089 (
            .in(out_3088),
            .outp(out_3089)
        );
        

        logic [WIDTH-1:0] out_3090;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3090 (
            .a(out_336),
            .b(out_3089),
            .outp(out_3090)
        );        
        

        logic [WIDTH-1:0] out_3091;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3091 (
            .a(out_3085),
            .b(out_3090),
            .outp(out_3091)
        );        
        

        logic [WIDTH-1:0] out_3092;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3092 (
            .a(out_3089),
            .b(out_343),
            .outp(out_3092)
        );        
        

        logic [WIDTH-1:0] out_3093;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3093 (
            .a(out_3091),
            .b(out_3092),
            .outp(out_3093)
        );        
        

        logic [WIDTH-1:0] out_3094;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3094 (
            .a(out_3093),
            .b(out_2892),
            .outp(out_3094)
        );        
        

        logic [WIDTH-1:0] out_3095;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3095 (
            .a(out_3083),
            .b(out_3094),
            .outp(out_3095)
        );        
        

        logic [WIDTH-1:0] out_3096;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.3)
        ) inst_3096 (
            .outp(out_3096)
        );
        

        logic [WIDTH-1:0] out_3097;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3097 (
            .a(out_14),
            .b(out_3096),
            .outp(out_3097)
        );        
        

        logic [WIDTH-1:0] out_3098;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.55)
        ) inst_3098 (
            .outp(out_3098)
        );
        

        logic [WIDTH-1:0] out_3099;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3099 (
            .a(out_3098),
            .b(out_14),
            .outp(out_3099)
        );        
        

        logic [WIDTH-1:0] out_3100;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3100 (
            .a(out_3097),
            .b(out_3099),
            .outp(out_3100)
        );        
        

        logic [WIDTH-1:0] out_3101;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.72551)
        ) inst_3101 (
            .outp(out_3101)
        );
        

        logic [WIDTH-1:0] out_3102;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3102 (
            .a(out_3),
            .b(out_3101),
            .outp(out_3102)
        );        
        

        logic [WIDTH-1:0] out_3103;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3103 (
            .a(out_3100),
            .b(out_3102),
            .outp(out_3103)
        );        
        

        logic [WIDTH-1:0] out_3104;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.62551)
        ) inst_3104 (
            .outp(out_3104)
        );
        

        logic [WIDTH-1:0] out_3105;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3105 (
            .a(out_3104),
            .b(out_3),
            .outp(out_3105)
        );        
        

        logic [WIDTH-1:0] out_3106;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3106 (
            .a(out_3103),
            .b(out_3105),
            .outp(out_3106)
        );        
        

        logic [WIDTH-1:0] out_3107;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3107 (
            .a(out_3095),
            .b(out_3106),
            .outp(out_3107)
        );        
        

        logic [WIDTH-1:0] out_3108;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.95)
        ) inst_3108 (
            .outp(out_3108)
        );
        

        logic [WIDTH-1:0] out_3109;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3109 (
            .a(out_14),
            .b(out_3108),
            .outp(out_3109)
        );        
        

        logic [WIDTH-1:0] out_3110;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.85)
        ) inst_3110 (
            .outp(out_3110)
        );
        

        logic [WIDTH-1:0] out_3111;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3111 (
            .a(out_3110),
            .b(out_14),
            .outp(out_3111)
        );        
        

        logic [WIDTH-1:0] out_3112;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3112 (
            .a(out_3109),
            .b(out_3111),
            .outp(out_3112)
        );        
        

        logic [WIDTH-1:0] out_3113;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.87551)
        ) inst_3113 (
            .outp(out_3113)
        );
        

        logic [WIDTH-1:0] out_3114;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3114 (
            .a(out_3),
            .b(out_3113),
            .outp(out_3114)
        );        
        

        logic [WIDTH-1:0] out_3115;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3115 (
            .a(out_3112),
            .b(out_3114),
            .outp(out_3115)
        );        
        

        logic [WIDTH-1:0] out_3116;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.47551)
        ) inst_3116 (
            .outp(out_3116)
        );
        

        logic [WIDTH-1:0] out_3117;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3117 (
            .a(out_3116),
            .b(out_3),
            .outp(out_3117)
        );        
        

        logic [WIDTH-1:0] out_3118;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3118 (
            .a(out_3115),
            .b(out_3117),
            .outp(out_3118)
        );        
        

        logic [WIDTH-1:0] out_3119;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3119 (
            .a(out_3107),
            .b(out_3118),
            .outp(out_3119)
        );        
        

        logic [WIDTH-1:0] out_3120;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3120 (
            .a(out_3114),
            .b(out_3117),
            .outp(out_3120)
        );        
        

        logic [WIDTH-1:0] out_3121;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3121 (
            .a(out_14),
            .b(out_3098),
            .outp(out_3121)
        );        
        

        logic [WIDTH-1:0] out_3122;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3122 (
            .a(out_3120),
            .b(out_3121),
            .outp(out_3122)
        );        
        

        logic [WIDTH-1:0] out_3123;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.3)
        ) inst_3123 (
            .outp(out_3123)
        );
        

        logic [WIDTH-1:0] out_3124;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3124 (
            .a(out_3123),
            .b(out_14),
            .outp(out_3124)
        );        
        

        logic [WIDTH-1:0] out_3125;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3125 (
            .a(out_3122),
            .b(out_3124),
            .outp(out_3125)
        );        
        

        logic [WIDTH-1:0] out_3126;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3126 (
            .in(out_3121),
            .outp(out_3126)
        );
        

        logic [WIDTH-1:0] out_3127;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3127 (
            .in(out_3114),
            .outp(out_3127)
        );
        

        logic [WIDTH-1:0] out_3128;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3128 (
            .a(out_3126),
            .b(out_3127),
            .outp(out_3128)
        );        
        

        logic [WIDTH-1:0] out_3129;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3129 (
            .in(out_3128),
            .outp(out_3129)
        );
        

        logic [WIDTH-1:0] out_3130;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3130 (
            .a(out_336),
            .b(out_3129),
            .outp(out_3130)
        );        
        

        logic [WIDTH-1:0] out_3131;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3131 (
            .a(out_3125),
            .b(out_3130),
            .outp(out_3131)
        );        
        

        logic [WIDTH-1:0] out_3132;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3132 (
            .a(out_3129),
            .b(out_343),
            .outp(out_3132)
        );        
        

        logic [WIDTH-1:0] out_3133;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3133 (
            .a(out_3131),
            .b(out_3132),
            .outp(out_3133)
        );        
        

        logic [WIDTH-1:0] out_3134;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3134 (
            .a(out_3119),
            .b(out_3133),
            .outp(out_3134)
        );        
        

        logic [WIDTH-1:0] out_3135;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.65)
        ) inst_3135 (
            .outp(out_3135)
        );
        

        logic [WIDTH-1:0] out_3136;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3136 (
            .a(out_14),
            .b(out_3135),
            .outp(out_3136)
        );        
        

        logic [WIDTH-1:0] out_3137;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3137 (
            .a(out_3124),
            .b(out_3136),
            .outp(out_3137)
        );        
        

        logic [WIDTH-1:0] out_3138;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.35551)
        ) inst_3138 (
            .outp(out_3138)
        );
        

        logic [WIDTH-1:0] out_3139;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3139 (
            .a(out_3),
            .b(out_3138),
            .outp(out_3139)
        );        
        

        logic [WIDTH-1:0] out_3140;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3140 (
            .a(out_3137),
            .b(out_3139),
            .outp(out_3140)
        );        
        

        logic [WIDTH-1:0] out_3141;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.25551)
        ) inst_3141 (
            .outp(out_3141)
        );
        

        logic [WIDTH-1:0] out_3142;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3142 (
            .a(out_3141),
            .b(out_3),
            .outp(out_3142)
        );        
        

        logic [WIDTH-1:0] out_3143;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3143 (
            .a(out_3140),
            .b(out_3142),
            .outp(out_3143)
        );        
        

        logic [WIDTH-1:0] out_3144;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3144 (
            .a(out_3134),
            .b(out_3143),
            .outp(out_3144)
        );        
        

        logic [WIDTH-1:0] out_3145;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.575)
        ) inst_3145 (
            .outp(out_3145)
        );
        

        logic [WIDTH-1:0] out_3146;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3146 (
            .a(out_14),
            .b(out_3145),
            .outp(out_3146)
        );        
        

        logic [WIDTH-1:0] out_3147;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3147 (
            .in(out_3146),
            .outp(out_3147)
        );
        

        logic [WIDTH-1:0] out_3148;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.90979)
        ) inst_3148 (
            .outp(out_3148)
        );
        

        logic [WIDTH-1:0] out_3149;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3149 (
            .a(out_1495),
            .b(out_3148),
            .outp(out_3149)
        );        
        

        logic [WIDTH-1:0] out_3150;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3150 (
            .a(out_3),
            .b(out_3149),
            .outp(out_3150)
        );        
        

        logic [WIDTH-1:0] out_3151;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3151 (
            .in(out_3150),
            .outp(out_3151)
        );
        

        logic [WIDTH-1:0] out_3152;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3152 (
            .a(out_3147),
            .b(out_3151),
            .outp(out_3152)
        );        
        

        logic [WIDTH-1:0] out_3153;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3153 (
            .in(out_3152),
            .outp(out_3153)
        );
        

        logic [WIDTH-1:0] out_3154;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3154 (
            .a(out_9),
            .b(out_3153),
            .outp(out_3154)
        );        
        

        logic [WIDTH-1:0] out_3155;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3155 (
            .a(out_3153),
            .b(out_21),
            .outp(out_3155)
        );        
        

        logic [WIDTH-1:0] out_3156;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3156 (
            .a(out_3154),
            .b(out_3155),
            .outp(out_3156)
        );        
        

        logic [WIDTH-1:0] out_3157;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3157 (
            .a(out_3144),
            .b(out_3156),
            .outp(out_3157)
        );        
        

        logic [WIDTH-1:0] out_3158;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.13393)
        ) inst_3158 (
            .outp(out_3158)
        );
        

        logic [WIDTH-1:0] out_3159;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3159 (
            .a(out_3158),
            .b(out_3),
            .outp(out_3159)
        );        
        

        logic [WIDTH-1:0] out_3160;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3160 (
            .a(out_3159),
            .b(out_1495),
            .outp(out_3160)
        );        
        

        logic [WIDTH-1:0] out_3161;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3161 (
            .in(out_3160),
            .outp(out_3161)
        );
        

        logic [WIDTH-1:0] out_3162;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3162 (
            .a(out_3161),
            .b(out_2962),
            .outp(out_3162)
        );        
        

        logic [WIDTH-1:0] out_3163;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3163 (
            .in(out_3162),
            .outp(out_3163)
        );
        

        logic [WIDTH-1:0] out_3164;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3164 (
            .a(out_9),
            .b(out_3163),
            .outp(out_3164)
        );        
        

        logic [WIDTH-1:0] out_3165;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3165 (
            .a(out_3163),
            .b(out_21),
            .outp(out_3165)
        );        
        

        logic [WIDTH-1:0] out_3166;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3166 (
            .a(out_3164),
            .b(out_3165),
            .outp(out_3166)
        );        
        

        logic [WIDTH-1:0] out_3167;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3167 (
            .a(out_3157),
            .b(out_3166),
            .outp(out_3167)
        );        
        

        logic [WIDTH-1:0] out_3168;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.7375)
        ) inst_3168 (
            .outp(out_3168)
        );
        

        logic [WIDTH-1:0] out_3169;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3169 (
            .a(out_3168),
            .b(out_260),
            .outp(out_3169)
        );        
        

        logic [WIDTH-1:0] out_3170;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3170 (
            .in(out_3169),
            .outp(out_3170)
        );
        

        logic [WIDTH-1:0] out_3171;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.575)
        ) inst_3171 (
            .outp(out_3171)
        );
        

        logic [WIDTH-1:0] out_3172;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3172 (
            .a(out_3171),
            .b(out_260),
            .outp(out_3172)
        );        
        

        logic [WIDTH-1:0] out_3173;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3173 (
            .a(out_3170),
            .b(out_3172),
            .outp(out_3173)
        );        
        

        logic [WIDTH-1:0] out_3174;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.575)
        ) inst_3174 (
            .outp(out_3174)
        );
        

        logic [WIDTH-1:0] out_3175;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3175 (
            .a(out_3174),
            .b(out_14),
            .outp(out_3175)
        );        
        

        logic [WIDTH-1:0] out_3176;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3176 (
            .in(out_3175),
            .outp(out_3176)
        );
        

        logic [WIDTH-1:0] out_3177;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3177 (
            .a(out_3173),
            .b(out_3176),
            .outp(out_3177)
        );        
        

        logic [WIDTH-1:0] out_3178;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4125)
        ) inst_3178 (
            .outp(out_3178)
        );
        

        logic [WIDTH-1:0] out_3179;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3179 (
            .a(out_3178),
            .b(out_14),
            .outp(out_3179)
        );        
        

        logic [WIDTH-1:0] out_3180;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3180 (
            .a(out_3177),
            .b(out_3179),
            .outp(out_3180)
        );        
        

        logic [WIDTH-1:0] out_3181;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.49333)
        ) inst_3181 (
            .outp(out_3181)
        );
        

        logic [WIDTH-1:0] out_3182;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3182 (
            .a(out_3181),
            .b(out_241),
            .outp(out_3182)
        );        
        

        logic [WIDTH-1:0] out_3183;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3183 (
            .in(out_3182),
            .outp(out_3183)
        );
        

        logic [WIDTH-1:0] out_3184;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3184 (
            .in(out_3183),
            .outp(out_3184)
        );
        

        logic [WIDTH-1:0] out_3185;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.415)
        ) inst_3185 (
            .outp(out_3185)
        );
        

        logic [WIDTH-1:0] out_3186;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3186 (
            .a(out_3185),
            .b(out_14),
            .outp(out_3186)
        );        
        

        logic [WIDTH-1:0] out_3187;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3187 (
            .in(out_3186),
            .outp(out_3187)
        );
        

        logic [WIDTH-1:0] out_3188;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3188 (
            .in(out_3187),
            .outp(out_3188)
        );
        

        logic [WIDTH-1:0] out_3189;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3189 (
            .a(out_3184),
            .b(out_3188),
            .outp(out_3189)
        );        
        

        logic [WIDTH-1:0] out_3190;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3190 (
            .in(out_3189),
            .outp(out_3190)
        );
        

        logic [WIDTH-1:0] out_3191;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3191 (
            .a(out_3190),
            .b(out_250),
            .outp(out_3191)
        );        
        

        logic [WIDTH-1:0] out_3192;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3192 (
            .a(out_3180),
            .b(out_3191),
            .outp(out_3192)
        );        
        

        logic [WIDTH-1:0] out_3193;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3193 (
            .in(out_3192),
            .outp(out_3193)
        );
        

        logic [WIDTH-1:0] out_3194;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3194 (
            .in(out_3170),
            .outp(out_3194)
        );
        

        logic [WIDTH-1:0] out_3195;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4125)
        ) inst_3195 (
            .outp(out_3195)
        );
        

        logic [WIDTH-1:0] out_3196;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3196 (
            .a(out_3195),
            .b(out_14),
            .outp(out_3196)
        );        
        

        logic [WIDTH-1:0] out_3197;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3197 (
            .in(out_3196),
            .outp(out_3197)
        );
        

        logic [WIDTH-1:0] out_3198;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3198 (
            .in(out_3197),
            .outp(out_3198)
        );
        

        logic [WIDTH-1:0] out_3199;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3199 (
            .a(out_3194),
            .b(out_3198),
            .outp(out_3199)
        );        
        

        logic [WIDTH-1:0] out_3200;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3200 (
            .in(out_3199),
            .outp(out_3200)
        );
        

        logic [WIDTH-1:0] out_3201;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3201 (
            .a(out_3200),
            .b(out_275),
            .outp(out_3201)
        );        
        

        logic [WIDTH-1:0] out_3202;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3202 (
            .a(out_3193),
            .b(out_3201),
            .outp(out_3202)
        );        
        

        logic [WIDTH-1:0] out_3203;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3203 (
            .a(out_3167),
            .b(out_3202),
            .outp(out_3203)
        );        
        

        logic [WIDTH-1:0] out_3204;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.7375)
        ) inst_3204 (
            .outp(out_3204)
        );
        

        logic [WIDTH-1:0] out_3205;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3205 (
            .a(out_3204),
            .b(out_260),
            .outp(out_3205)
        );        
        

        logic [WIDTH-1:0] out_3206;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.9)
        ) inst_3206 (
            .outp(out_3206)
        );
        

        logic [WIDTH-1:0] out_3207;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3207 (
            .a(out_3206),
            .b(out_260),
            .outp(out_3207)
        );        
        

        logic [WIDTH-1:0] out_3208;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3208 (
            .in(out_3207),
            .outp(out_3208)
        );
        

        logic [WIDTH-1:0] out_3209;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3209 (
            .a(out_3205),
            .b(out_3208),
            .outp(out_3209)
        );        
        

        logic [WIDTH-1:0] out_3210;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.475)
        ) inst_3210 (
            .outp(out_3210)
        );
        

        logic [WIDTH-1:0] out_3211;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3211 (
            .a(out_3210),
            .b(out_14),
            .outp(out_3211)
        );        
        

        logic [WIDTH-1:0] out_3212;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3212 (
            .a(out_3209),
            .b(out_3211),
            .outp(out_3212)
        );        
        

        logic [WIDTH-1:0] out_3213;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6375)
        ) inst_3213 (
            .outp(out_3213)
        );
        

        logic [WIDTH-1:0] out_3214;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3214 (
            .a(out_3213),
            .b(out_14),
            .outp(out_3214)
        );        
        

        logic [WIDTH-1:0] out_3215;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3215 (
            .in(out_3214),
            .outp(out_3215)
        );
        

        logic [WIDTH-1:0] out_3216;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3216 (
            .a(out_3212),
            .b(out_3215),
            .outp(out_3216)
        );        
        

        logic [WIDTH-1:0] out_3217;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.49)
        ) inst_3217 (
            .outp(out_3217)
        );
        

        logic [WIDTH-1:0] out_3218;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3218 (
            .a(out_3217),
            .b(out_241),
            .outp(out_3218)
        );        
        

        logic [WIDTH-1:0] out_3219;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3219 (
            .in(out_3218),
            .outp(out_3219)
        );
        

        logic [WIDTH-1:0] out_3220;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.635)
        ) inst_3220 (
            .outp(out_3220)
        );
        

        logic [WIDTH-1:0] out_3221;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3221 (
            .a(out_3220),
            .b(out_14),
            .outp(out_3221)
        );        
        

        logic [WIDTH-1:0] out_3222;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3222 (
            .in(out_3221),
            .outp(out_3222)
        );
        

        logic [WIDTH-1:0] out_3223;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3223 (
            .a(out_3219),
            .b(out_3222),
            .outp(out_3223)
        );        
        

        logic [WIDTH-1:0] out_3224;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3224 (
            .in(out_3223),
            .outp(out_3224)
        );
        

        logic [WIDTH-1:0] out_3225;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3225 (
            .a(out_3224),
            .b(out_250),
            .outp(out_3225)
        );        
        

        logic [WIDTH-1:0] out_3226;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3226 (
            .a(out_3216),
            .b(out_3225),
            .outp(out_3226)
        );        
        

        logic [WIDTH-1:0] out_3227;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3227 (
            .in(out_3226),
            .outp(out_3227)
        );
        

        logic [WIDTH-1:0] out_3228;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3228 (
            .in(out_3205),
            .outp(out_3228)
        );
        

        logic [WIDTH-1:0] out_3229;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6375)
        ) inst_3229 (
            .outp(out_3229)
        );
        

        logic [WIDTH-1:0] out_3230;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3230 (
            .a(out_3229),
            .b(out_14),
            .outp(out_3230)
        );        
        

        logic [WIDTH-1:0] out_3231;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3231 (
            .in(out_3230),
            .outp(out_3231)
        );
        

        logic [WIDTH-1:0] out_3232;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3232 (
            .a(out_3228),
            .b(out_3231),
            .outp(out_3232)
        );        
        

        logic [WIDTH-1:0] out_3233;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3233 (
            .in(out_3232),
            .outp(out_3233)
        );
        

        logic [WIDTH-1:0] out_3234;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3234 (
            .a(out_3233),
            .b(out_275),
            .outp(out_3234)
        );        
        

        logic [WIDTH-1:0] out_3235;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3235 (
            .a(out_3227),
            .b(out_3234),
            .outp(out_3235)
        );        
        

        logic [WIDTH-1:0] out_3236;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3236 (
            .a(out_3203),
            .b(out_3235),
            .outp(out_3236)
        );        
        

        logic [WIDTH-1:0] out_3237;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.075)
        ) inst_3237 (
            .outp(out_3237)
        );
        

        logic [WIDTH-1:0] out_3238;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3238 (
            .a(out_3237),
            .b(out_3),
            .outp(out_3238)
        );        
        

        logic [WIDTH-1:0] out_3239;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3239 (
            .in(out_3238),
            .outp(out_3239)
        );
        

        logic [WIDTH-1:0] out_3240;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.975)
        ) inst_3240 (
            .outp(out_3240)
        );
        

        logic [WIDTH-1:0] out_3241;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3241 (
            .a(out_3240),
            .b(out_3),
            .outp(out_3241)
        );        
        

        logic [WIDTH-1:0] out_3242;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3242 (
            .a(out_3239),
            .b(out_3241),
            .outp(out_3242)
        );        
        

        logic [WIDTH-1:0] out_3243;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3243 (
            .a(out_3242),
            .b(out_2888),
            .outp(out_3243)
        );        
        

        logic [WIDTH-1:0] out_3244;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3244 (
            .a(out_3243),
            .b(out_2892),
            .outp(out_3244)
        );        
        

        logic [WIDTH-1:0] out_3245;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3245 (
            .a(out_3236),
            .b(out_3244),
            .outp(out_3245)
        );        
        

        logic [WIDTH-1:0] out_3246;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.025)
        ) inst_3246 (
            .outp(out_3246)
        );
        

        logic [WIDTH-1:0] out_3247;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3247 (
            .a(out_3246),
            .b(out_3),
            .outp(out_3247)
        );        
        

        logic [WIDTH-1:0] out_3248;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3248 (
            .in(out_3247),
            .outp(out_3248)
        );
        

        logic [WIDTH-1:0] out_3249;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3249 (
            .a(out_3248),
            .b(out_2931),
            .outp(out_3249)
        );        
        

        logic [WIDTH-1:0] out_3250;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3250 (
            .in(out_3249),
            .outp(out_3250)
        );
        

        logic [WIDTH-1:0] out_3251;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3251 (
            .a(out_3250),
            .b(out_460),
            .outp(out_3251)
        );        
        

        logic [WIDTH-1:0] out_3252;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3252 (
            .a(out_3245),
            .b(out_3251),
            .outp(out_3252)
        );        
        

        logic [WIDTH-1:0] out_3253;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.35)
        ) inst_3253 (
            .outp(out_3253)
        );
        

        logic [WIDTH-1:0] out_3254;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3254 (
            .a(out_3253),
            .b(out_3),
            .outp(out_3254)
        );        
        

        logic [WIDTH-1:0] out_3255;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3255 (
            .in(out_3254),
            .outp(out_3255)
        );
        

        logic [WIDTH-1:0] out_3256;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3256 (
            .a(out_3041),
            .b(out_3255),
            .outp(out_3256)
        );        
        

        logic [WIDTH-1:0] out_3257;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3257 (
            .a(out_3256),
            .b(out_2961),
            .outp(out_3257)
        );        
        

        logic [WIDTH-1:0] out_3258;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3258 (
            .a(out_3257),
            .b(out_2892),
            .outp(out_3258)
        );        
        

        logic [WIDTH-1:0] out_3259;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3259 (
            .a(out_3252),
            .b(out_3258),
            .outp(out_3259)
        );        
        

        logic [WIDTH-1:0] out_3260;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.7)
        ) inst_3260 (
            .outp(out_3260)
        );
        

        logic [WIDTH-1:0] out_3261;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3261 (
            .a(out_3260),
            .b(out_3),
            .outp(out_3261)
        );        
        

        logic [WIDTH-1:0] out_3262;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3262 (
            .a(out_3261),
            .b(out_3045),
            .outp(out_3262)
        );        
        

        logic [WIDTH-1:0] out_3263;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3263 (
            .a(out_3262),
            .b(out_2985),
            .outp(out_3263)
        );        
        

        logic [WIDTH-1:0] out_3264;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3264 (
            .a(out_3263),
            .b(out_2892),
            .outp(out_3264)
        );        
        

        logic [WIDTH-1:0] out_3265;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3265 (
            .a(out_3259),
            .b(out_3264),
            .outp(out_3265)
        );        
        

        logic [WIDTH-1:0] out_3266;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3266 (
            .a(out_14),
            .b(out_669),
            .outp(out_3266)
        );        
        

        logic [WIDTH-1:0] out_3267;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3267 (
            .in(out_3266),
            .outp(out_3267)
        );
        

        logic [WIDTH-1:0] out_3268;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.02467)
        ) inst_3268 (
            .outp(out_3268)
        );
        

        logic [WIDTH-1:0] out_3269;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3269 (
            .a(out_241),
            .b(out_3268),
            .outp(out_3269)
        );        
        

        logic [WIDTH-1:0] out_3270;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3270 (
            .in(out_3269),
            .outp(out_3270)
        );
        

        logic [WIDTH-1:0] out_3271;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3271 (
            .a(out_3267),
            .b(out_3270),
            .outp(out_3271)
        );        
        

        logic [WIDTH-1:0] out_3272;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3272 (
            .in(out_3271),
            .outp(out_3272)
        );
        

        logic [WIDTH-1:0] out_3273;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3273 (
            .a(out_3272),
            .b(out_250),
            .outp(out_3273)
        );        
        

        logic [WIDTH-1:0] out_3274;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.625)
        ) inst_3274 (
            .outp(out_3274)
        );
        

        logic [WIDTH-1:0] out_3275;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3275 (
            .a(out_14),
            .b(out_3274),
            .outp(out_3275)
        );        
        

        logic [WIDTH-1:0] out_3276;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4625)
        ) inst_3276 (
            .outp(out_3276)
        );
        

        logic [WIDTH-1:0] out_3277;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3277 (
            .a(out_3276),
            .b(out_14),
            .outp(out_3277)
        );        
        

        logic [WIDTH-1:0] out_3278;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3278 (
            .a(out_3275),
            .b(out_3277),
            .outp(out_3278)
        );        
        

        logic [WIDTH-1:0] out_3279;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0345)
        ) inst_3279 (
            .outp(out_3279)
        );
        

        logic [WIDTH-1:0] out_3280;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3280 (
            .a(out_260),
            .b(out_3279),
            .outp(out_3280)
        );        
        

        logic [WIDTH-1:0] out_3281;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3281 (
            .a(out_3278),
            .b(out_3280),
            .outp(out_3281)
        );        
        

        logic [WIDTH-1:0] out_3282;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.872)
        ) inst_3282 (
            .outp(out_3282)
        );
        

        logic [WIDTH-1:0] out_3283;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3283 (
            .a(out_3282),
            .b(out_260),
            .outp(out_3283)
        );        
        

        logic [WIDTH-1:0] out_3284;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3284 (
            .a(out_3281),
            .b(out_3283),
            .outp(out_3284)
        );        
        

        logic [WIDTH-1:0] out_3285;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3285 (
            .a(out_3273),
            .b(out_3284),
            .outp(out_3285)
        );        
        

        logic [WIDTH-1:0] out_3286;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3286 (
            .in(out_3285),
            .outp(out_3286)
        );
        

        logic [WIDTH-1:0] out_3287;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4625)
        ) inst_3287 (
            .outp(out_3287)
        );
        

        logic [WIDTH-1:0] out_3288;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3288 (
            .a(out_14),
            .b(out_3287),
            .outp(out_3288)
        );        
        

        logic [WIDTH-1:0] out_3289;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3289 (
            .in(out_3288),
            .outp(out_3289)
        );
        

        logic [WIDTH-1:0] out_3290;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3290 (
            .in(out_3280),
            .outp(out_3290)
        );
        

        logic [WIDTH-1:0] out_3291;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3291 (
            .a(out_3289),
            .b(out_3290),
            .outp(out_3291)
        );        
        

        logic [WIDTH-1:0] out_3292;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3292 (
            .in(out_3291),
            .outp(out_3292)
        );
        

        logic [WIDTH-1:0] out_3293;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3293 (
            .a(out_3292),
            .b(out_275),
            .outp(out_3293)
        );        
        

        logic [WIDTH-1:0] out_3294;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3294 (
            .a(out_3286),
            .b(out_3293),
            .outp(out_3294)
        );        
        

        logic [WIDTH-1:0] out_3295;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3295 (
            .a(out_3265),
            .b(out_3294),
            .outp(out_3295)
        );        
        

        logic [WIDTH-1:0] out_3296;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.615)
        ) inst_3296 (
            .outp(out_3296)
        );
        

        logic [WIDTH-1:0] out_3297;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3297 (
            .a(out_14),
            .b(out_3296),
            .outp(out_3297)
        );        
        

        logic [WIDTH-1:0] out_3298;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.525)
        ) inst_3298 (
            .outp(out_3298)
        );
        

        logic [WIDTH-1:0] out_3299;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3299 (
            .a(out_3298),
            .b(out_14),
            .outp(out_3299)
        );        
        

        logic [WIDTH-1:0] out_3300;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3300 (
            .a(out_3297),
            .b(out_3299),
            .outp(out_3300)
        );        
        

        logic [WIDTH-1:0] out_3301;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.208)
        ) inst_3301 (
            .outp(out_3301)
        );
        

        logic [WIDTH-1:0] out_3302;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3302 (
            .a(out_3),
            .b(out_3301),
            .outp(out_3302)
        );        
        

        logic [WIDTH-1:0] out_3303;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3303 (
            .a(out_3300),
            .b(out_3302),
            .outp(out_3303)
        );        
        

        logic [WIDTH-1:0] out_3304;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.708)
        ) inst_3304 (
            .outp(out_3304)
        );
        

        logic [WIDTH-1:0] out_3305;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3305 (
            .a(out_3304),
            .b(out_3),
            .outp(out_3305)
        );        
        

        logic [WIDTH-1:0] out_3306;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3306 (
            .a(out_3303),
            .b(out_3305),
            .outp(out_3306)
        );        
        

        logic [WIDTH-1:0] out_3307;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.933)
        ) inst_3307 (
            .outp(out_3307)
        );
        

        logic [WIDTH-1:0] out_3308;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3308 (
            .a(out_3),
            .b(out_3307),
            .outp(out_3308)
        );        
        

        logic [WIDTH-1:0] out_3309;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3309 (
            .in(out_3308),
            .outp(out_3309)
        );
        

        logic [WIDTH-1:0] out_3310;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3310 (
            .a(out_3147),
            .b(out_3309),
            .outp(out_3310)
        );        
        

        logic [WIDTH-1:0] out_3311;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3311 (
            .in(out_3310),
            .outp(out_3311)
        );
        

        logic [WIDTH-1:0] out_3312;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3312 (
            .a(out_3311),
            .b(out_21),
            .outp(out_3312)
        );        
        

        logic [WIDTH-1:0] out_3313;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.37375)
        ) inst_3313 (
            .outp(out_3313)
        );
        

        logic [WIDTH-1:0] out_3314;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3314 (
            .a(out_553),
            .b(out_3313),
            .outp(out_3314)
        );        
        

        logic [WIDTH-1:0] out_3315;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.12595)
        ) inst_3315 (
            .outp(out_3315)
        );
        

        logic [WIDTH-1:0] out_3316;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3316 (
            .a(out_3315),
            .b(out_559),
            .outp(out_3316)
        );        
        

        logic [WIDTH-1:0] out_3317;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3317 (
            .a(out_556),
            .b(out_3316),
            .outp(out_3317)
        );        
        

        logic [WIDTH-1:0] out_3318;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3318 (
            .a(out_3314),
            .b(out_3317),
            .outp(out_3318)
        );        
        

        logic [WIDTH-1:0] out_3319;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.32095)
        ) inst_3319 (
            .outp(out_3319)
        );
        

        logic [WIDTH-1:0] out_3320;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3320 (
            .a(out_3319),
            .b(out_2653),
            .outp(out_3320)
        );        
        

        logic [WIDTH-1:0] out_3321;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3321 (
            .a(out_3318),
            .b(out_3320),
            .outp(out_3321)
        );        
        

        logic [WIDTH-1:0] out_3322;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3322 (
            .a(out_2653),
            .b(out_3319),
            .outp(out_3322)
        );        
        

        logic [WIDTH-1:0] out_3323;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3323 (
            .a(out_3316),
            .b(out_556),
            .outp(out_3323)
        );        
        

        logic [WIDTH-1:0] out_3324;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3324 (
            .a(out_3322),
            .b(out_3323),
            .outp(out_3324)
        );        
        

        logic [WIDTH-1:0] out_3325;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3325 (
            .a(out_3313),
            .b(out_553),
            .outp(out_3325)
        );        
        

        logic [WIDTH-1:0] out_3326;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3326 (
            .a(out_3324),
            .b(out_3325),
            .outp(out_3326)
        );        
        

        logic [WIDTH-1:0] out_3327;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3327 (
            .a(out_3321),
            .b(out_3326),
            .outp(out_3327)
        );        
        

        logic [WIDTH-1:0] out_3328;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3328 (
            .in(out_3327),
            .outp(out_3328)
        );
        

        logic [WIDTH-1:0] out_3329;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3329 (
            .a(out_3312),
            .b(out_3328),
            .outp(out_3329)
        );        
        

        logic [WIDTH-1:0] out_3330;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3330 (
            .a(out_9),
            .b(out_3311),
            .outp(out_3330)
        );        
        

        logic [WIDTH-1:0] out_3331;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3331 (
            .a(out_3329),
            .b(out_3330),
            .outp(out_3331)
        );        
        

        logic [WIDTH-1:0] out_3332;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3332 (
            .a(out_3306),
            .b(out_3331),
            .outp(out_3332)
        );        
        

        logic [WIDTH-1:0] out_3333;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3333 (
            .a(out_3312),
            .b(out_3332),
            .outp(out_3333)
        );        
        

        logic [WIDTH-1:0] out_3334;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3334 (
            .a(out_3295),
            .b(out_3333),
            .outp(out_3334)
        );        
        

        logic [WIDTH-1:0] out_3335;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.2095)
        ) inst_3335 (
            .outp(out_3335)
        );
        

        logic [WIDTH-1:0] out_3336;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3336 (
            .a(out_3335),
            .b(out_260),
            .outp(out_3336)
        );        
        

        logic [WIDTH-1:0] out_3337;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.372)
        ) inst_3337 (
            .outp(out_3337)
        );
        

        logic [WIDTH-1:0] out_3338;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3338 (
            .a(out_260),
            .b(out_3337),
            .outp(out_3338)
        );        
        

        logic [WIDTH-1:0] out_3339;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3339 (
            .a(out_3336),
            .b(out_3338),
            .outp(out_3339)
        );        
        

        logic [WIDTH-1:0] out_3340;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.525)
        ) inst_3340 (
            .outp(out_3340)
        );
        

        logic [WIDTH-1:0] out_3341;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3341 (
            .a(out_3340),
            .b(out_14),
            .outp(out_3341)
        );        
        

        logic [WIDTH-1:0] out_3342;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3342 (
            .a(out_3339),
            .b(out_3341),
            .outp(out_3342)
        );        
        

        logic [WIDTH-1:0] out_3343;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6875)
        ) inst_3343 (
            .outp(out_3343)
        );
        

        logic [WIDTH-1:0] out_3344;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3344 (
            .a(out_14),
            .b(out_3343),
            .outp(out_3344)
        );        
        

        logic [WIDTH-1:0] out_3345;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3345 (
            .a(out_3342),
            .b(out_3344),
            .outp(out_3345)
        );        
        

        logic [WIDTH-1:0] out_3346;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.47133)
        ) inst_3346 (
            .outp(out_3346)
        );
        

        logic [WIDTH-1:0] out_3347;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3347 (
            .a(out_3346),
            .b(out_241),
            .outp(out_3347)
        );        
        

        logic [WIDTH-1:0] out_3348;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3348 (
            .in(out_3347),
            .outp(out_3348)
        );
        

        logic [WIDTH-1:0] out_3349;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.685)
        ) inst_3349 (
            .outp(out_3349)
        );
        

        logic [WIDTH-1:0] out_3350;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3350 (
            .a(out_3349),
            .b(out_14),
            .outp(out_3350)
        );        
        

        logic [WIDTH-1:0] out_3351;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3351 (
            .in(out_3350),
            .outp(out_3351)
        );
        

        logic [WIDTH-1:0] out_3352;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3352 (
            .a(out_3348),
            .b(out_3351),
            .outp(out_3352)
        );        
        

        logic [WIDTH-1:0] out_3353;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3353 (
            .in(out_3352),
            .outp(out_3353)
        );
        

        logic [WIDTH-1:0] out_3354;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3354 (
            .a(out_3353),
            .b(out_250),
            .outp(out_3354)
        );        
        

        logic [WIDTH-1:0] out_3355;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3355 (
            .a(out_3345),
            .b(out_3354),
            .outp(out_3355)
        );        
        

        logic [WIDTH-1:0] out_3356;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3356 (
            .in(out_3355),
            .outp(out_3356)
        );
        

        logic [WIDTH-1:0] out_3357;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3357 (
            .in(out_3336),
            .outp(out_3357)
        );
        

        logic [WIDTH-1:0] out_3358;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6875)
        ) inst_3358 (
            .outp(out_3358)
        );
        

        logic [WIDTH-1:0] out_3359;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3359 (
            .a(out_3358),
            .b(out_14),
            .outp(out_3359)
        );        
        

        logic [WIDTH-1:0] out_3360;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3360 (
            .in(out_3359),
            .outp(out_3360)
        );
        

        logic [WIDTH-1:0] out_3361;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3361 (
            .a(out_3357),
            .b(out_3360),
            .outp(out_3361)
        );        
        

        logic [WIDTH-1:0] out_3362;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3362 (
            .in(out_3361),
            .outp(out_3362)
        );
        

        logic [WIDTH-1:0] out_3363;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3363 (
            .a(out_3362),
            .b(out_275),
            .outp(out_3363)
        );        
        

        logic [WIDTH-1:0] out_3364;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3364 (
            .a(out_3356),
            .b(out_3363),
            .outp(out_3364)
        );        
        

        logic [WIDTH-1:0] out_3365;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3365 (
            .a(out_3334),
            .b(out_3364),
            .outp(out_3365)
        );        
        

        logic [WIDTH-1:0] out_3366;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3366 (
            .a(out_3124),
            .b(out_3146),
            .outp(out_3366)
        );        
        

        logic [WIDTH-1:0] out_3367;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.6455)
        ) inst_3367 (
            .outp(out_3367)
        );
        

        logic [WIDTH-1:0] out_3368;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3368 (
            .a(out_3),
            .b(out_3367),
            .outp(out_3368)
        );        
        

        logic [WIDTH-1:0] out_3369;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3369 (
            .a(out_3366),
            .b(out_3368),
            .outp(out_3369)
        );        
        

        logic [WIDTH-1:0] out_3370;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.5455)
        ) inst_3370 (
            .outp(out_3370)
        );
        

        logic [WIDTH-1:0] out_3371;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3371 (
            .a(out_3370),
            .b(out_3),
            .outp(out_3371)
        );        
        

        logic [WIDTH-1:0] out_3372;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3372 (
            .a(out_3369),
            .b(out_3371),
            .outp(out_3372)
        );        
        

        logic [WIDTH-1:0] out_3373;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3373 (
            .a(out_3365),
            .b(out_3372),
            .outp(out_3373)
        );        
        

        logic [WIDTH-1:0] out_3374;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3374 (
            .a(out_3097),
            .b(out_3124),
            .outp(out_3374)
        );        
        

        logic [WIDTH-1:0] out_3375;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.19551)
        ) inst_3375 (
            .outp(out_3375)
        );
        

        logic [WIDTH-1:0] out_3376;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3376 (
            .a(out_3),
            .b(out_3375),
            .outp(out_3376)
        );        
        

        logic [WIDTH-1:0] out_3377;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3377 (
            .a(out_3374),
            .b(out_3376),
            .outp(out_3377)
        );        
        

        logic [WIDTH-1:0] out_3378;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.0955)
        ) inst_3378 (
            .outp(out_3378)
        );
        

        logic [WIDTH-1:0] out_3379;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3379 (
            .a(out_3378),
            .b(out_3),
            .outp(out_3379)
        );        
        

        logic [WIDTH-1:0] out_3380;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3380 (
            .a(out_3377),
            .b(out_3379),
            .outp(out_3380)
        );        
        

        logic [WIDTH-1:0] out_3381;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3381 (
            .a(out_3373),
            .b(out_3380),
            .outp(out_3381)
        );        
        

        logic [WIDTH-1:0] out_3382;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3382 (
            .a(out_3368),
            .b(out_3379),
            .outp(out_3382)
        );        
        

        logic [WIDTH-1:0] out_3383;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.85)
        ) inst_3383 (
            .outp(out_3383)
        );
        

        logic [WIDTH-1:0] out_3384;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3384 (
            .a(out_14),
            .b(out_3383),
            .outp(out_3384)
        );        
        

        logic [WIDTH-1:0] out_3385;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3385 (
            .a(out_3382),
            .b(out_3384),
            .outp(out_3385)
        );        
        

        logic [WIDTH-1:0] out_3386;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3386 (
            .a(out_135),
            .b(out_14),
            .outp(out_3386)
        );        
        

        logic [WIDTH-1:0] out_3387;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3387 (
            .a(out_3385),
            .b(out_3386),
            .outp(out_3387)
        );        
        

        logic [WIDTH-1:0] out_3388;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.3705)
        ) inst_3388 (
            .outp(out_3388)
        );
        

        logic [WIDTH-1:0] out_3389;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3389 (
            .a(out_3),
            .b(out_3388),
            .outp(out_3389)
        );        
        

        logic [WIDTH-1:0] out_3390;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3390 (
            .in(out_3389),
            .outp(out_3390)
        );
        

        logic [WIDTH-1:0] out_3391;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3391 (
            .a(out_3147),
            .b(out_3390),
            .outp(out_3391)
        );        
        

        logic [WIDTH-1:0] out_3392;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3392 (
            .in(out_3391),
            .outp(out_3392)
        );
        

        logic [WIDTH-1:0] out_3393;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3393 (
            .a(out_9),
            .b(out_3392),
            .outp(out_3393)
        );        
        

        logic [WIDTH-1:0] out_3394;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3394 (
            .a(out_3387),
            .b(out_3393),
            .outp(out_3394)
        );        
        

        logic [WIDTH-1:0] out_3395;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3395 (
            .a(out_3392),
            .b(out_21),
            .outp(out_3395)
        );        
        

        logic [WIDTH-1:0] out_3396;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3396 (
            .a(out_3394),
            .b(out_3395),
            .outp(out_3396)
        );        
        

        logic [WIDTH-1:0] out_3397;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3397 (
            .a(out_3381),
            .b(out_3396),
            .outp(out_3397)
        );        
        

        logic [WIDTH-1:0] out_3398;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.8455)
        ) inst_3398 (
            .outp(out_3398)
        );
        

        logic [WIDTH-1:0] out_3399;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3399 (
            .a(out_3),
            .b(out_3398),
            .outp(out_3399)
        );        
        

        logic [WIDTH-1:0] out_3400;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3400 (
            .a(out_3100),
            .b(out_3399),
            .outp(out_3400)
        );        
        

        logic [WIDTH-1:0] out_3401;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.7455)
        ) inst_3401 (
            .outp(out_3401)
        );
        

        logic [WIDTH-1:0] out_3402;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3402 (
            .a(out_3401),
            .b(out_3),
            .outp(out_3402)
        );        
        

        logic [WIDTH-1:0] out_3403;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3403 (
            .a(out_3400),
            .b(out_3402),
            .outp(out_3403)
        );        
        

        logic [WIDTH-1:0] out_3404;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3404 (
            .a(out_3397),
            .b(out_3403),
            .outp(out_3404)
        );        
        

        logic [WIDTH-1:0] out_3405;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.9955)
        ) inst_3405 (
            .outp(out_3405)
        );
        

        logic [WIDTH-1:0] out_3406;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3406 (
            .a(out_3),
            .b(out_3405),
            .outp(out_3406)
        );        
        

        logic [WIDTH-1:0] out_3407;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3407 (
            .a(out_3112),
            .b(out_3406),
            .outp(out_3407)
        );        
        

        logic [WIDTH-1:0] out_3408;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.5955)
        ) inst_3408 (
            .outp(out_3408)
        );
        

        logic [WIDTH-1:0] out_3409;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3409 (
            .a(out_3408),
            .b(out_3),
            .outp(out_3409)
        );        
        

        logic [WIDTH-1:0] out_3410;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3410 (
            .a(out_3407),
            .b(out_3409),
            .outp(out_3410)
        );        
        

        logic [WIDTH-1:0] out_3411;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3411 (
            .a(out_3404),
            .b(out_3410),
            .outp(out_3411)
        );        
        

        logic [WIDTH-1:0] out_3412;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3412 (
            .a(out_3121),
            .b(out_3124),
            .outp(out_3412)
        );        
        

        logic [WIDTH-1:0] out_3413;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3413 (
            .a(out_3412),
            .b(out_3406),
            .outp(out_3413)
        );        
        

        logic [WIDTH-1:0] out_3414;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3414 (
            .a(out_3413),
            .b(out_3409),
            .outp(out_3414)
        );        
        

        logic [WIDTH-1:0] out_3415;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3415 (
            .in(out_3406),
            .outp(out_3415)
        );
        

        logic [WIDTH-1:0] out_3416;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3416 (
            .a(out_3126),
            .b(out_3415),
            .outp(out_3416)
        );        
        

        logic [WIDTH-1:0] out_3417;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3417 (
            .in(out_3416),
            .outp(out_3417)
        );
        

        logic [WIDTH-1:0] out_3418;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3418 (
            .a(out_336),
            .b(out_3417),
            .outp(out_3418)
        );        
        

        logic [WIDTH-1:0] out_3419;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3419 (
            .a(out_3414),
            .b(out_3418),
            .outp(out_3419)
        );        
        

        logic [WIDTH-1:0] out_3420;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3420 (
            .a(out_3417),
            .b(out_343),
            .outp(out_3420)
        );        
        

        logic [WIDTH-1:0] out_3421;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3421 (
            .a(out_3419),
            .b(out_3420),
            .outp(out_3421)
        );        
        

        logic [WIDTH-1:0] out_3422;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3422 (
            .a(out_3411),
            .b(out_3421),
            .outp(out_3422)
        );        
        

        logic [WIDTH-1:0] out_3423;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3423 (
            .a(out_3341),
            .b(out_3344),
            .outp(out_3423)
        );        
        

        logic [WIDTH-1:0] out_3424;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0345)
        ) inst_3424 (
            .outp(out_3424)
        );
        

        logic [WIDTH-1:0] out_3425;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3425 (
            .a(out_3424),
            .b(out_260),
            .outp(out_3425)
        );        
        

        logic [WIDTH-1:0] out_3426;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3426 (
            .a(out_3423),
            .b(out_3425),
            .outp(out_3426)
        );        
        

        logic [WIDTH-1:0] out_3427;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.197)
        ) inst_3427 (
            .outp(out_3427)
        );
        

        logic [WIDTH-1:0] out_3428;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3428 (
            .a(out_260),
            .b(out_3427),
            .outp(out_3428)
        );        
        

        logic [WIDTH-1:0] out_3429;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3429 (
            .a(out_3426),
            .b(out_3428),
            .outp(out_3429)
        );        
        

        logic [WIDTH-1:0] out_3430;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.02133)
        ) inst_3430 (
            .outp(out_3430)
        );
        

        logic [WIDTH-1:0] out_3431;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3431 (
            .a(out_3430),
            .b(out_241),
            .outp(out_3431)
        );        
        

        logic [WIDTH-1:0] out_3432;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3432 (
            .in(out_3431),
            .outp(out_3432)
        );
        

        logic [WIDTH-1:0] out_3433;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3433 (
            .a(out_3351),
            .b(out_3432),
            .outp(out_3433)
        );        
        

        logic [WIDTH-1:0] out_3434;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3434 (
            .in(out_3433),
            .outp(out_3434)
        );
        

        logic [WIDTH-1:0] out_3435;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3435 (
            .a(out_3434),
            .b(out_250),
            .outp(out_3435)
        );        
        

        logic [WIDTH-1:0] out_3436;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3436 (
            .a(out_3429),
            .b(out_3435),
            .outp(out_3436)
        );        
        

        logic [WIDTH-1:0] out_3437;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3437 (
            .in(out_3436),
            .outp(out_3437)
        );
        

        logic [WIDTH-1:0] out_3438;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3438 (
            .in(out_3425),
            .outp(out_3438)
        );
        

        logic [WIDTH-1:0] out_3439;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3439 (
            .a(out_3360),
            .b(out_3438),
            .outp(out_3439)
        );        
        

        logic [WIDTH-1:0] out_3440;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3440 (
            .in(out_3439),
            .outp(out_3440)
        );
        

        logic [WIDTH-1:0] out_3441;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3441 (
            .a(out_3440),
            .b(out_275),
            .outp(out_3441)
        );        
        

        logic [WIDTH-1:0] out_3442;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3442 (
            .a(out_3437),
            .b(out_3441),
            .outp(out_3442)
        );        
        

        logic [WIDTH-1:0] out_3443;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3443 (
            .a(out_3422),
            .b(out_3442),
            .outp(out_3443)
        );        
        

        logic [WIDTH-1:0] out_3444;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.788667)
        ) inst_3444 (
            .outp(out_3444)
        );
        

        logic [WIDTH-1:0] out_3445;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3445 (
            .a(out_3444),
            .b(out_260),
            .outp(out_3445)
        );        
        

        logic [WIDTH-1:0] out_3446;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3446 (
            .a(out_3278),
            .b(out_3445),
            .outp(out_3446)
        );        
        

        logic [WIDTH-1:0] out_3447;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.951167)
        ) inst_3447 (
            .outp(out_3447)
        );
        

        logic [WIDTH-1:0] out_3448;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3448 (
            .a(out_260),
            .b(out_3447),
            .outp(out_3448)
        );        
        

        logic [WIDTH-1:0] out_3449;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3449 (
            .a(out_3446),
            .b(out_3448),
            .outp(out_3449)
        );        
        

        logic [WIDTH-1:0] out_3450;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.635778)
        ) inst_3450 (
            .outp(out_3450)
        );
        

        logic [WIDTH-1:0] out_3451;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3451 (
            .a(out_241),
            .b(out_3450),
            .outp(out_3451)
        );        
        

        logic [WIDTH-1:0] out_3452;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3452 (
            .in(out_3451),
            .outp(out_3452)
        );
        

        logic [WIDTH-1:0] out_3453;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3453 (
            .a(out_3267),
            .b(out_3452),
            .outp(out_3453)
        );        
        

        logic [WIDTH-1:0] out_3454;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3454 (
            .in(out_3453),
            .outp(out_3454)
        );
        

        logic [WIDTH-1:0] out_3455;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3455 (
            .a(out_3454),
            .b(out_250),
            .outp(out_3455)
        );        
        

        logic [WIDTH-1:0] out_3456;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3456 (
            .a(out_3449),
            .b(out_3455),
            .outp(out_3456)
        );        
        

        logic [WIDTH-1:0] out_3457;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3457 (
            .in(out_3456),
            .outp(out_3457)
        );
        

        logic [WIDTH-1:0] out_3458;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3458 (
            .in(out_3448),
            .outp(out_3458)
        );
        

        logic [WIDTH-1:0] out_3459;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3459 (
            .a(out_3289),
            .b(out_3458),
            .outp(out_3459)
        );        
        

        logic [WIDTH-1:0] out_3460;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3460 (
            .in(out_3459),
            .outp(out_3460)
        );
        

        logic [WIDTH-1:0] out_3461;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3461 (
            .a(out_3460),
            .b(out_275),
            .outp(out_3461)
        );        
        

        logic [WIDTH-1:0] out_3462;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3462 (
            .a(out_3457),
            .b(out_3461),
            .outp(out_3462)
        );        
        

        logic [WIDTH-1:0] out_3463;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3463 (
            .a(out_3443),
            .b(out_3462),
            .outp(out_3463)
        );        
        

        logic [WIDTH-1:0] out_3464;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3464 (
            .a(out_3124),
            .b(out_3384),
            .outp(out_3464)
        );        
        

        logic [WIDTH-1:0] out_3465;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.125)
        ) inst_3465 (
            .outp(out_3465)
        );
        

        logic [WIDTH-1:0] out_3466;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3466 (
            .a(out_3),
            .b(out_3465),
            .outp(out_3466)
        );        
        

        logic [WIDTH-1:0] out_3467;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3467 (
            .a(out_3464),
            .b(out_3466),
            .outp(out_3467)
        );        
        

        logic [WIDTH-1:0] out_3468;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0249996)
        ) inst_3468 (
            .outp(out_3468)
        );
        

        logic [WIDTH-1:0] out_3469;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3469 (
            .a(out_3468),
            .b(out_3),
            .outp(out_3469)
        );        
        

        logic [WIDTH-1:0] out_3470;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3470 (
            .a(out_3467),
            .b(out_3469),
            .outp(out_3470)
        );        
        

        logic [WIDTH-1:0] out_3471;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3471 (
            .a(out_3463),
            .b(out_3470),
            .outp(out_3471)
        );        
        

        logic [WIDTH-1:0] out_3472;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.585714)
        ) inst_3472 (
            .outp(out_3472)
        );
        

        logic [WIDTH-1:0] out_3473;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3473 (
            .a(out_194),
            .b(out_3472),
            .outp(out_3473)
        );        
        

        logic [WIDTH-1:0] out_3474;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3474 (
            .a(out_3464),
            .b(out_3473),
            .outp(out_3474)
        );        
        

        logic [WIDTH-1:0] out_3475;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0357141)
        ) inst_3475 (
            .outp(out_3475)
        );
        

        logic [WIDTH-1:0] out_3476;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3476 (
            .a(out_3475),
            .b(out_194),
            .outp(out_3476)
        );        
        

        logic [WIDTH-1:0] out_3477;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3477 (
            .a(out_3474),
            .b(out_3476),
            .outp(out_3477)
        );        
        

        logic [WIDTH-1:0] out_3478;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3478 (
            .a(out_14),
            .b(out_3123),
            .outp(out_3478)
        );        
        

        logic [WIDTH-1:0] out_3479;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3479 (
            .in(out_3478),
            .outp(out_3479)
        );
        

        logic [WIDTH-1:0] out_3480;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.732143)
        ) inst_3480 (
            .outp(out_3480)
        );
        

        logic [WIDTH-1:0] out_3481;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3481 (
            .a(out_204),
            .b(out_3480),
            .outp(out_3481)
        );        
        

        logic [WIDTH-1:0] out_3482;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3482 (
            .in(out_3481),
            .outp(out_3482)
        );
        

        logic [WIDTH-1:0] out_3483;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3483 (
            .a(out_3479),
            .b(out_3482),
            .outp(out_3483)
        );        
        

        logic [WIDTH-1:0] out_3484;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3484 (
            .in(out_3483),
            .outp(out_3484)
        );
        

        logic [WIDTH-1:0] out_3485;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3485 (
            .a(out_200),
            .b(out_3484),
            .outp(out_3485)
        );        
        

        logic [WIDTH-1:0] out_3486;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3486 (
            .a(out_3477),
            .b(out_3485),
            .outp(out_3486)
        );        
        

        logic [WIDTH-1:0] out_3487;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3487 (
            .in(out_3473),
            .outp(out_3487)
        );
        

        logic [WIDTH-1:0] out_3488;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3488 (
            .a(out_3479),
            .b(out_3487),
            .outp(out_3488)
        );        
        

        logic [WIDTH-1:0] out_3489;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3489 (
            .in(out_3488),
            .outp(out_3489)
        );
        

        logic [WIDTH-1:0] out_3490;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3490 (
            .a(out_3489),
            .b(out_214),
            .outp(out_3490)
        );        
        

        logic [WIDTH-1:0] out_3491;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3491 (
            .a(out_3486),
            .b(out_3490),
            .outp(out_3491)
        );        
        

        logic [WIDTH-1:0] out_3492;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3492 (
            .a(out_3471),
            .b(out_3491),
            .outp(out_3492)
        );        
        

        logic [WIDTH-1:0] out_3493;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.1)
        ) inst_3493 (
            .outp(out_3493)
        );
        

        logic [WIDTH-1:0] out_3494;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3494 (
            .a(out_3493),
            .b(out_3),
            .outp(out_3494)
        );        
        

        logic [WIDTH-1:0] out_3495;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3495 (
            .a(out_3464),
            .b(out_3494),
            .outp(out_3495)
        );        
        

        logic [WIDTH-1:0] out_3496;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.2)
        ) inst_3496 (
            .outp(out_3496)
        );
        

        logic [WIDTH-1:0] out_3497;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3497 (
            .a(out_3496),
            .b(out_3),
            .outp(out_3497)
        );        
        

        logic [WIDTH-1:0] out_3498;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3498 (
            .in(out_3497),
            .outp(out_3498)
        );
        

        logic [WIDTH-1:0] out_3499;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3499 (
            .a(out_3495),
            .b(out_3498),
            .outp(out_3499)
        );        
        

        logic [WIDTH-1:0] out_3500;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3500 (
            .a(out_3492),
            .b(out_3499),
            .outp(out_3500)
        );        
        

        logic [WIDTH-1:0] out_3501;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.0)
        ) inst_3501 (
            .outp(out_3501)
        );
        

        logic [WIDTH-1:0] out_3502;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3502 (
            .a(out_14),
            .b(out_3501),
            .outp(out_3502)
        );        
        

        logic [WIDTH-1:0] out_3503;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3503 (
            .in(out_3502),
            .outp(out_3503)
        );
        

        logic [WIDTH-1:0] out_3504;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.150001)
        ) inst_3504 (
            .outp(out_3504)
        );
        

        logic [WIDTH-1:0] out_3505;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3505 (
            .a(out_3504),
            .b(out_3),
            .outp(out_3505)
        );        
        

        logic [WIDTH-1:0] out_3506;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3506 (
            .in(out_3505),
            .outp(out_3506)
        );
        

        logic [WIDTH-1:0] out_3507;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3507 (
            .a(out_3503),
            .b(out_3506),
            .outp(out_3507)
        );        
        

        logic [WIDTH-1:0] out_3508;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3508 (
            .in(out_3507),
            .outp(out_3508)
        );
        

        logic [WIDTH-1:0] out_3509;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3509 (
            .a(out_3508),
            .b(out_460),
            .outp(out_3509)
        );        
        

        logic [WIDTH-1:0] out_3510;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3510 (
            .a(out_3500),
            .b(out_3509),
            .outp(out_3510)
        );        
        

        logic [WIDTH-1:0] out_3511;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.325)
        ) inst_3511 (
            .outp(out_3511)
        );
        

        logic [WIDTH-1:0] out_3512;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3512 (
            .a(out_3511),
            .b(out_3),
            .outp(out_3512)
        );        
        

        logic [WIDTH-1:0] out_3513;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3513 (
            .a(out_3300),
            .b(out_3512),
            .outp(out_3513)
        );        
        

        logic [WIDTH-1:0] out_3514;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.825)
        ) inst_3514 (
            .outp(out_3514)
        );
        

        logic [WIDTH-1:0] out_3515;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3515 (
            .a(out_3514),
            .b(out_3),
            .outp(out_3515)
        );        
        

        logic [WIDTH-1:0] out_3516;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3516 (
            .in(out_3515),
            .outp(out_3516)
        );
        

        logic [WIDTH-1:0] out_3517;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3517 (
            .a(out_3513),
            .b(out_3516),
            .outp(out_3517)
        );        
        

        logic [WIDTH-1:0] out_3518;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6)
        ) inst_3518 (
            .outp(out_3518)
        );
        

        logic [WIDTH-1:0] out_3519;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3519 (
            .a(out_3518),
            .b(out_3),
            .outp(out_3519)
        );        
        

        logic [WIDTH-1:0] out_3520;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3520 (
            .in(out_3519),
            .outp(out_3520)
        );
        

        logic [WIDTH-1:0] out_3521;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3521 (
            .a(out_3147),
            .b(out_3520),
            .outp(out_3521)
        );        
        

        logic [WIDTH-1:0] out_3522;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3522 (
            .in(out_3521),
            .outp(out_3522)
        );
        

        logic [WIDTH-1:0] out_3523;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3523 (
            .a(out_3522),
            .b(out_21),
            .outp(out_3523)
        );        
        

        logic [WIDTH-1:0] out_3524;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.120625)
        ) inst_3524 (
            .outp(out_3524)
        );
        

        logic [WIDTH-1:0] out_3525;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3525 (
            .a(out_3524),
            .b(out_556),
            .outp(out_3525)
        );        
        

        logic [WIDTH-1:0] out_3526;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3526 (
            .a(out_3525),
            .b(out_559),
            .outp(out_3526)
        );        
        

        logic [WIDTH-1:0] out_3527;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3527 (
            .a(out_3314),
            .b(out_3526),
            .outp(out_3527)
        );        
        

        logic [WIDTH-1:0] out_3528;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0743749)
        ) inst_3528 (
            .outp(out_3528)
        );
        

        logic [WIDTH-1:0] out_3529;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3529 (
            .a(out_3528),
            .b(out_2653),
            .outp(out_3529)
        );        
        

        logic [WIDTH-1:0] out_3530;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3530 (
            .a(out_3527),
            .b(out_3529),
            .outp(out_3530)
        );        
        

        logic [WIDTH-1:0] out_3531;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3531 (
            .a(out_2653),
            .b(out_3528),
            .outp(out_3531)
        );        
        

        logic [WIDTH-1:0] out_3532;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3532 (
            .a(out_3325),
            .b(out_3531),
            .outp(out_3532)
        );        
        

        logic [WIDTH-1:0] out_3533;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3533 (
            .a(out_559),
            .b(out_3525),
            .outp(out_3533)
        );        
        

        logic [WIDTH-1:0] out_3534;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3534 (
            .a(out_3532),
            .b(out_3533),
            .outp(out_3534)
        );        
        

        logic [WIDTH-1:0] out_3535;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3535 (
            .a(out_3530),
            .b(out_3534),
            .outp(out_3535)
        );        
        

        logic [WIDTH-1:0] out_3536;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3536 (
            .in(out_3535),
            .outp(out_3536)
        );
        

        logic [WIDTH-1:0] out_3537;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3537 (
            .a(out_3523),
            .b(out_3536),
            .outp(out_3537)
        );        
        

        logic [WIDTH-1:0] out_3538;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3538 (
            .a(out_9),
            .b(out_3522),
            .outp(out_3538)
        );        
        

        logic [WIDTH-1:0] out_3539;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3539 (
            .a(out_3537),
            .b(out_3538),
            .outp(out_3539)
        );        
        

        logic [WIDTH-1:0] out_3540;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3540 (
            .a(out_3517),
            .b(out_3539),
            .outp(out_3540)
        );        
        

        logic [WIDTH-1:0] out_3541;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3541 (
            .a(out_3523),
            .b(out_3540),
            .outp(out_3541)
        );        
        

        logic [WIDTH-1:0] out_3542;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3542 (
            .a(out_3510),
            .b(out_3541),
            .outp(out_3542)
        );        
        

        logic [WIDTH-1:0] out_3543;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.2095)
        ) inst_3543 (
            .outp(out_3543)
        );
        

        logic [WIDTH-1:0] out_3544;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3544 (
            .a(out_260),
            .b(out_3543),
            .outp(out_3544)
        );        
        

        logic [WIDTH-1:0] out_3545;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.047)
        ) inst_3545 (
            .outp(out_3545)
        );
        

        logic [WIDTH-1:0] out_3546;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3546 (
            .a(out_3545),
            .b(out_260),
            .outp(out_3546)
        );        
        

        logic [WIDTH-1:0] out_3547;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3547 (
            .a(out_3544),
            .b(out_3546),
            .outp(out_3547)
        );        
        

        logic [WIDTH-1:0] out_3548;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3548 (
            .a(out_3547),
            .b(out_3275),
            .outp(out_3548)
        );        
        

        logic [WIDTH-1:0] out_3549;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3549 (
            .a(out_3548),
            .b(out_3277),
            .outp(out_3549)
        );        
        

        logic [WIDTH-1:0] out_3550;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.47467)
        ) inst_3550 (
            .outp(out_3550)
        );
        

        logic [WIDTH-1:0] out_3551;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3551 (
            .a(out_241),
            .b(out_3550),
            .outp(out_3551)
        );        
        

        logic [WIDTH-1:0] out_3552;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3552 (
            .in(out_3551),
            .outp(out_3552)
        );
        

        logic [WIDTH-1:0] out_3553;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3553 (
            .a(out_3267),
            .b(out_3552),
            .outp(out_3553)
        );        
        

        logic [WIDTH-1:0] out_3554;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3554 (
            .in(out_3553),
            .outp(out_3554)
        );
        

        logic [WIDTH-1:0] out_3555;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3555 (
            .a(out_3554),
            .b(out_250),
            .outp(out_3555)
        );        
        

        logic [WIDTH-1:0] out_3556;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3556 (
            .a(out_3549),
            .b(out_3555),
            .outp(out_3556)
        );        
        

        logic [WIDTH-1:0] out_3557;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3557 (
            .in(out_3556),
            .outp(out_3557)
        );
        

        logic [WIDTH-1:0] out_3558;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3558 (
            .in(out_3544),
            .outp(out_3558)
        );
        

        logic [WIDTH-1:0] out_3559;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3559 (
            .a(out_3289),
            .b(out_3558),
            .outp(out_3559)
        );        
        

        logic [WIDTH-1:0] out_3560;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3560 (
            .in(out_3559),
            .outp(out_3560)
        );
        

        logic [WIDTH-1:0] out_3561;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3561 (
            .a(out_3560),
            .b(out_275),
            .outp(out_3561)
        );        
        

        logic [WIDTH-1:0] out_3562;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3562 (
            .a(out_3557),
            .b(out_3561),
            .outp(out_3562)
        );        
        

        logic [WIDTH-1:0] out_3563;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3563 (
            .a(out_3542),
            .b(out_3562),
            .outp(out_3563)
        );        
        

        logic [WIDTH-1:0] out_3564;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3564 (
            .a(out_3124),
            .b(out_3275),
            .outp(out_3564)
        );        
        

        logic [WIDTH-1:0] out_3565;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.9705)
        ) inst_3565 (
            .outp(out_3565)
        );
        

        logic [WIDTH-1:0] out_3566;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3566 (
            .a(out_3),
            .b(out_3565),
            .outp(out_3566)
        );        
        

        logic [WIDTH-1:0] out_3567;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3567 (
            .a(out_3564),
            .b(out_3566),
            .outp(out_3567)
        );        
        

        logic [WIDTH-1:0] out_3568;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8705)
        ) inst_3568 (
            .outp(out_3568)
        );
        

        logic [WIDTH-1:0] out_3569;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3569 (
            .a(out_3568),
            .b(out_3),
            .outp(out_3569)
        );        
        

        logic [WIDTH-1:0] out_3570;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3570 (
            .a(out_3567),
            .b(out_3569),
            .outp(out_3570)
        );        
        

        logic [WIDTH-1:0] out_3571;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3571 (
            .a(out_3563),
            .b(out_3570),
            .outp(out_3571)
        );        
        

        logic [WIDTH-1:0] out_3572;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5205)
        ) inst_3572 (
            .outp(out_3572)
        );
        

        logic [WIDTH-1:0] out_3573;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3573 (
            .a(out_3),
            .b(out_3572),
            .outp(out_3573)
        );        
        

        logic [WIDTH-1:0] out_3574;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3574 (
            .a(out_3464),
            .b(out_3573),
            .outp(out_3574)
        );        
        

        logic [WIDTH-1:0] out_3575;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.4205)
        ) inst_3575 (
            .outp(out_3575)
        );
        

        logic [WIDTH-1:0] out_3576;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3576 (
            .a(out_3575),
            .b(out_3),
            .outp(out_3576)
        );        
        

        logic [WIDTH-1:0] out_3577;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3577 (
            .a(out_3574),
            .b(out_3576),
            .outp(out_3577)
        );        
        

        logic [WIDTH-1:0] out_3578;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3578 (
            .a(out_3571),
            .b(out_3577),
            .outp(out_3578)
        );        
        

        logic [WIDTH-1:0] out_3579;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3579 (
            .a(out_3384),
            .b(out_3566),
            .outp(out_3579)
        );        
        

        logic [WIDTH-1:0] out_3580;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3580 (
            .a(out_3579),
            .b(out_3576),
            .outp(out_3580)
        );        
        

        logic [WIDTH-1:0] out_3581;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.625)
        ) inst_3581 (
            .outp(out_3581)
        );
        

        logic [WIDTH-1:0] out_3582;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3582 (
            .a(out_3581),
            .b(out_14),
            .outp(out_3582)
        );        
        

        logic [WIDTH-1:0] out_3583;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3583 (
            .a(out_3580),
            .b(out_3582),
            .outp(out_3583)
        );        
        

        logic [WIDTH-1:0] out_3584;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6955)
        ) inst_3584 (
            .outp(out_3584)
        );
        

        logic [WIDTH-1:0] out_3585;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3585 (
            .a(out_3),
            .b(out_3584),
            .outp(out_3585)
        );        
        

        logic [WIDTH-1:0] out_3586;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3586 (
            .in(out_3585),
            .outp(out_3586)
        );
        

        logic [WIDTH-1:0] out_3587;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3587 (
            .a(out_3147),
            .b(out_3586),
            .outp(out_3587)
        );        
        

        logic [WIDTH-1:0] out_3588;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3588 (
            .in(out_3587),
            .outp(out_3588)
        );
        

        logic [WIDTH-1:0] out_3589;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3589 (
            .a(out_9),
            .b(out_3588),
            .outp(out_3589)
        );        
        

        logic [WIDTH-1:0] out_3590;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3590 (
            .a(out_3583),
            .b(out_3589),
            .outp(out_3590)
        );        
        

        logic [WIDTH-1:0] out_3591;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3591 (
            .a(out_3588),
            .b(out_21),
            .outp(out_3591)
        );        
        

        logic [WIDTH-1:0] out_3592;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3592 (
            .a(out_3590),
            .b(out_3591),
            .outp(out_3592)
        );        
        

        logic [WIDTH-1:0] out_3593;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3593 (
            .a(out_3578),
            .b(out_3592),
            .outp(out_3593)
        );        
        

        logic [WIDTH-1:0] out_3594;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.3205)
        ) inst_3594 (
            .outp(out_3594)
        );
        

        logic [WIDTH-1:0] out_3595;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3595 (
            .a(out_3),
            .b(out_3594),
            .outp(out_3595)
        );        
        

        logic [WIDTH-1:0] out_3596;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3596 (
            .a(out_3300),
            .b(out_3595),
            .outp(out_3596)
        );        
        

        logic [WIDTH-1:0] out_3597;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.8205)
        ) inst_3597 (
            .outp(out_3597)
        );
        

        logic [WIDTH-1:0] out_3598;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3598 (
            .a(out_3597),
            .b(out_3),
            .outp(out_3598)
        );        
        

        logic [WIDTH-1:0] out_3599;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3599 (
            .a(out_3596),
            .b(out_3598),
            .outp(out_3599)
        );        
        

        logic [WIDTH-1:0] out_3600;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0455)
        ) inst_3600 (
            .outp(out_3600)
        );
        

        logic [WIDTH-1:0] out_3601;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3601 (
            .a(out_3),
            .b(out_3600),
            .outp(out_3601)
        );        
        

        logic [WIDTH-1:0] out_3602;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3602 (
            .in(out_3601),
            .outp(out_3602)
        );
        

        logic [WIDTH-1:0] out_3603;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3603 (
            .a(out_3147),
            .b(out_3602),
            .outp(out_3603)
        );        
        

        logic [WIDTH-1:0] out_3604;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3604 (
            .in(out_3603),
            .outp(out_3604)
        );
        

        logic [WIDTH-1:0] out_3605;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3605 (
            .a(out_3604),
            .b(out_21),
            .outp(out_3605)
        );        
        

        logic [WIDTH-1:0] out_3606;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.606888)
        ) inst_3606 (
            .outp(out_3606)
        );
        

        logic [WIDTH-1:0] out_3607;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3607 (
            .a(out_3606),
            .b(out_559),
            .outp(out_3607)
        );        
        

        logic [WIDTH-1:0] out_3608;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3608 (
            .a(out_556),
            .b(out_3607),
            .outp(out_3608)
        );        
        

        logic [WIDTH-1:0] out_3609;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3609 (
            .a(out_3314),
            .b(out_3608),
            .outp(out_3609)
        );        
        

        logic [WIDTH-1:0] out_3610;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.801888)
        ) inst_3610 (
            .outp(out_3610)
        );
        

        logic [WIDTH-1:0] out_3611;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3611 (
            .a(out_3610),
            .b(out_2653),
            .outp(out_3611)
        );        
        

        logic [WIDTH-1:0] out_3612;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3612 (
            .a(out_3609),
            .b(out_3611),
            .outp(out_3612)
        );        
        

        logic [WIDTH-1:0] out_3613;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3613 (
            .a(out_2653),
            .b(out_3610),
            .outp(out_3613)
        );        
        

        logic [WIDTH-1:0] out_3614;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3614 (
            .a(out_3325),
            .b(out_3613),
            .outp(out_3614)
        );        
        

        logic [WIDTH-1:0] out_3615;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.606888)
        ) inst_3615 (
            .outp(out_3615)
        );
        

        logic [WIDTH-1:0] out_3616;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3616 (
            .a(out_3615),
            .b(out_559),
            .outp(out_3616)
        );        
        

        logic [WIDTH-1:0] out_3617;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3617 (
            .a(out_3616),
            .b(out_556),
            .outp(out_3617)
        );        
        

        logic [WIDTH-1:0] out_3618;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3618 (
            .a(out_3614),
            .b(out_3617),
            .outp(out_3618)
        );        
        

        logic [WIDTH-1:0] out_3619;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3619 (
            .a(out_3612),
            .b(out_3618),
            .outp(out_3619)
        );        
        

        logic [WIDTH-1:0] out_3620;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3620 (
            .in(out_3619),
            .outp(out_3620)
        );
        

        logic [WIDTH-1:0] out_3621;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3621 (
            .a(out_3605),
            .b(out_3620),
            .outp(out_3621)
        );        
        

        logic [WIDTH-1:0] out_3622;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3622 (
            .a(out_9),
            .b(out_3604),
            .outp(out_3622)
        );        
        

        logic [WIDTH-1:0] out_3623;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3623 (
            .a(out_3621),
            .b(out_3622),
            .outp(out_3623)
        );        
        

        logic [WIDTH-1:0] out_3624;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3624 (
            .a(out_3599),
            .b(out_3623),
            .outp(out_3624)
        );        
        

        logic [WIDTH-1:0] out_3625;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3625 (
            .a(out_3605),
            .b(out_3624),
            .outp(out_3625)
        );        
        

        logic [WIDTH-1:0] out_3626;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3626 (
            .a(out_3593),
            .b(out_3625),
            .outp(out_3626)
        );        
        

        logic [WIDTH-1:0] out_3627;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.951167)
        ) inst_3627 (
            .outp(out_3627)
        );
        

        logic [WIDTH-1:0] out_3628;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3628 (
            .a(out_3627),
            .b(out_260),
            .outp(out_3628)
        );        
        

        logic [WIDTH-1:0] out_3629;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3629 (
            .a(out_3423),
            .b(out_3628),
            .outp(out_3629)
        );        
        

        logic [WIDTH-1:0] out_3630;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.11367)
        ) inst_3630 (
            .outp(out_3630)
        );
        

        logic [WIDTH-1:0] out_3631;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3631 (
            .a(out_260),
            .b(out_3630),
            .outp(out_3631)
        );        
        

        logic [WIDTH-1:0] out_3632;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3632 (
            .a(out_3629),
            .b(out_3631),
            .outp(out_3632)
        );        
        

        logic [WIDTH-1:0] out_3633;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.632445)
        ) inst_3633 (
            .outp(out_3633)
        );
        

        logic [WIDTH-1:0] out_3634;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3634 (
            .a(out_3633),
            .b(out_241),
            .outp(out_3634)
        );        
        

        logic [WIDTH-1:0] out_3635;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3635 (
            .in(out_3634),
            .outp(out_3635)
        );
        

        logic [WIDTH-1:0] out_3636;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3636 (
            .a(out_3351),
            .b(out_3635),
            .outp(out_3636)
        );        
        

        logic [WIDTH-1:0] out_3637;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3637 (
            .in(out_3636),
            .outp(out_3637)
        );
        

        logic [WIDTH-1:0] out_3638;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3638 (
            .a(out_3637),
            .b(out_250),
            .outp(out_3638)
        );        
        

        logic [WIDTH-1:0] out_3639;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3639 (
            .a(out_3632),
            .b(out_3638),
            .outp(out_3639)
        );        
        

        logic [WIDTH-1:0] out_3640;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3640 (
            .in(out_3639),
            .outp(out_3640)
        );
        

        logic [WIDTH-1:0] out_3641;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3641 (
            .in(out_3628),
            .outp(out_3641)
        );
        

        logic [WIDTH-1:0] out_3642;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3642 (
            .a(out_3360),
            .b(out_3641),
            .outp(out_3642)
        );        
        

        logic [WIDTH-1:0] out_3643;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3643 (
            .in(out_3642),
            .outp(out_3643)
        );
        

        logic [WIDTH-1:0] out_3644;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3644 (
            .a(out_3643),
            .b(out_275),
            .outp(out_3644)
        );        
        

        logic [WIDTH-1:0] out_3645;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3645 (
            .a(out_3640),
            .b(out_3644),
            .outp(out_3645)
        );        
        

        logic [WIDTH-1:0] out_3646;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3646 (
            .a(out_3626),
            .b(out_3645),
            .outp(out_3646)
        );        
        

        logic [WIDTH-1:0] out_3647;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5125)
        ) inst_3647 (
            .outp(out_3647)
        );
        

        logic [WIDTH-1:0] out_3648;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3648 (
            .a(out_3647),
            .b(out_14),
            .outp(out_3648)
        );        
        

        logic [WIDTH-1:0] out_3649;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3649 (
            .in(out_3648),
            .outp(out_3649)
        );
        

        logic [WIDTH-1:0] out_3650;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3650 (
            .in(out_3649),
            .outp(out_3650)
        );
        

        logic [WIDTH-1:0] out_3651;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.3955)
        ) inst_3651 (
            .outp(out_3651)
        );
        

        logic [WIDTH-1:0] out_3652;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3652 (
            .a(out_3651),
            .b(out_260),
            .outp(out_3652)
        );        
        

        logic [WIDTH-1:0] out_3653;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3653 (
            .in(out_3652),
            .outp(out_3653)
        );
        

        logic [WIDTH-1:0] out_3654;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3654 (
            .in(out_3653),
            .outp(out_3654)
        );
        

        logic [WIDTH-1:0] out_3655;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3655 (
            .a(out_3650),
            .b(out_3654),
            .outp(out_3655)
        );        
        

        logic [WIDTH-1:0] out_3656;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3656 (
            .in(out_3655),
            .outp(out_3656)
        );
        

        logic [WIDTH-1:0] out_3657;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3657 (
            .a(out_3656),
            .b(out_275),
            .outp(out_3657)
        );        
        

        logic [WIDTH-1:0] out_3658;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.675)
        ) inst_3658 (
            .outp(out_3658)
        );
        

        logic [WIDTH-1:0] out_3659;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3659 (
            .a(out_3658),
            .b(out_14),
            .outp(out_3659)
        );        
        

        logic [WIDTH-1:0] out_3660;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3660 (
            .in(out_3659),
            .outp(out_3660)
        );
        

        logic [WIDTH-1:0] out_3661;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5125)
        ) inst_3661 (
            .outp(out_3661)
        );
        

        logic [WIDTH-1:0] out_3662;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3662 (
            .a(out_3661),
            .b(out_14),
            .outp(out_3662)
        );        
        

        logic [WIDTH-1:0] out_3663;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3663 (
            .a(out_3660),
            .b(out_3662),
            .outp(out_3663)
        );        
        

        logic [WIDTH-1:0] out_3664;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3664 (
            .a(out_3663),
            .b(out_3653),
            .outp(out_3664)
        );        
        

        logic [WIDTH-1:0] out_3665;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.233001)
        ) inst_3665 (
            .outp(out_3665)
        );
        

        logic [WIDTH-1:0] out_3666;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3666 (
            .a(out_3665),
            .b(out_260),
            .outp(out_3666)
        );        
        

        logic [WIDTH-1:0] out_3667;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3667 (
            .a(out_3664),
            .b(out_3666),
            .outp(out_3667)
        );        
        

        logic [WIDTH-1:0] out_3668;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.515)
        ) inst_3668 (
            .outp(out_3668)
        );
        

        logic [WIDTH-1:0] out_3669;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3669 (
            .a(out_3668),
            .b(out_14),
            .outp(out_3669)
        );        
        

        logic [WIDTH-1:0] out_3670;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3670 (
            .in(out_3669),
            .outp(out_3670)
        );
        

        logic [WIDTH-1:0] out_3671;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3671 (
            .in(out_3670),
            .outp(out_3671)
        );
        

        logic [WIDTH-1:0] out_3672;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.265334)
        ) inst_3672 (
            .outp(out_3672)
        );
        

        logic [WIDTH-1:0] out_3673;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3673 (
            .a(out_3672),
            .b(out_241),
            .outp(out_3673)
        );        
        

        logic [WIDTH-1:0] out_3674;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3674 (
            .in(out_3673),
            .outp(out_3674)
        );
        

        logic [WIDTH-1:0] out_3675;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3675 (
            .in(out_3674),
            .outp(out_3675)
        );
        

        logic [WIDTH-1:0] out_3676;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3676 (
            .a(out_3671),
            .b(out_3675),
            .outp(out_3676)
        );        
        

        logic [WIDTH-1:0] out_3677;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3677 (
            .in(out_3676),
            .outp(out_3677)
        );
        

        logic [WIDTH-1:0] out_3678;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3678 (
            .a(out_3677),
            .b(out_250),
            .outp(out_3678)
        );        
        

        logic [WIDTH-1:0] out_3679;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3679 (
            .a(out_3667),
            .b(out_3678),
            .outp(out_3679)
        );        
        

        logic [WIDTH-1:0] out_3680;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3680 (
            .in(out_3679),
            .outp(out_3680)
        );
        

        logic [WIDTH-1:0] out_3681;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3681 (
            .a(out_3657),
            .b(out_3680),
            .outp(out_3681)
        );        
        

        logic [WIDTH-1:0] out_3682;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3682 (
            .a(out_3646),
            .b(out_3681),
            .outp(out_3682)
        );        
        

        logic [WIDTH-1:0] out_3683;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.575)
        ) inst_3683 (
            .outp(out_3683)
        );
        

        logic [WIDTH-1:0] out_3684;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3684 (
            .a(out_3683),
            .b(out_14),
            .outp(out_3684)
        );        
        

        logic [WIDTH-1:0] out_3685;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.7375)
        ) inst_3685 (
            .outp(out_3685)
        );
        

        logic [WIDTH-1:0] out_3686;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3686 (
            .a(out_3685),
            .b(out_14),
            .outp(out_3686)
        );        
        

        logic [WIDTH-1:0] out_3687;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3687 (
            .in(out_3686),
            .outp(out_3687)
        );
        

        logic [WIDTH-1:0] out_3688;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3688 (
            .a(out_3684),
            .b(out_3687),
            .outp(out_3688)
        );        
        

        logic [WIDTH-1:0] out_3689;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.395501)
        ) inst_3689 (
            .outp(out_3689)
        );
        

        logic [WIDTH-1:0] out_3690;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3690 (
            .a(out_3689),
            .b(out_260),
            .outp(out_3690)
        );        
        

        logic [WIDTH-1:0] out_3691;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3691 (
            .a(out_3688),
            .b(out_3690),
            .outp(out_3691)
        );        
        

        logic [WIDTH-1:0] out_3692;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3692 (
            .a(out_593),
            .b(out_260),
            .outp(out_3692)
        );        
        

        logic [WIDTH-1:0] out_3693;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3693 (
            .in(out_3692),
            .outp(out_3693)
        );
        

        logic [WIDTH-1:0] out_3694;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3694 (
            .a(out_3691),
            .b(out_3693),
            .outp(out_3694)
        );        
        

        logic [WIDTH-1:0] out_3695;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.735)
        ) inst_3695 (
            .outp(out_3695)
        );
        

        logic [WIDTH-1:0] out_3696;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3696 (
            .a(out_3695),
            .b(out_14),
            .outp(out_3696)
        );        
        

        logic [WIDTH-1:0] out_3697;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3697 (
            .in(out_3696),
            .outp(out_3697)
        );
        

        logic [WIDTH-1:0] out_3698;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.262)
        ) inst_3698 (
            .outp(out_3698)
        );
        

        logic [WIDTH-1:0] out_3699;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3699 (
            .a(out_3698),
            .b(out_241),
            .outp(out_3699)
        );        
        

        logic [WIDTH-1:0] out_3700;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3700 (
            .in(out_3699),
            .outp(out_3700)
        );
        

        logic [WIDTH-1:0] out_3701;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3701 (
            .a(out_3697),
            .b(out_3700),
            .outp(out_3701)
        );        
        

        logic [WIDTH-1:0] out_3702;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3702 (
            .in(out_3701),
            .outp(out_3702)
        );
        

        logic [WIDTH-1:0] out_3703;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3703 (
            .a(out_3702),
            .b(out_250),
            .outp(out_3703)
        );        
        

        logic [WIDTH-1:0] out_3704;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3704 (
            .a(out_3694),
            .b(out_3703),
            .outp(out_3704)
        );        
        

        logic [WIDTH-1:0] out_3705;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3705 (
            .in(out_3704),
            .outp(out_3705)
        );
        

        logic [WIDTH-1:0] out_3706;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.7375)
        ) inst_3706 (
            .outp(out_3706)
        );
        

        logic [WIDTH-1:0] out_3707;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3707 (
            .a(out_3706),
            .b(out_14),
            .outp(out_3707)
        );        
        

        logic [WIDTH-1:0] out_3708;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3708 (
            .in(out_3707),
            .outp(out_3708)
        );
        

        logic [WIDTH-1:0] out_3709;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3709 (
            .in(out_3690),
            .outp(out_3709)
        );
        

        logic [WIDTH-1:0] out_3710;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3710 (
            .a(out_3708),
            .b(out_3709),
            .outp(out_3710)
        );        
        

        logic [WIDTH-1:0] out_3711;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3711 (
            .in(out_3710),
            .outp(out_3711)
        );
        

        logic [WIDTH-1:0] out_3712;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3712 (
            .a(out_3711),
            .b(out_275),
            .outp(out_3712)
        );        
        

        logic [WIDTH-1:0] out_3713;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3713 (
            .a(out_3705),
            .b(out_3712),
            .outp(out_3713)
        );        
        

        logic [WIDTH-1:0] out_3714;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3714 (
            .a(out_3682),
            .b(out_3713),
            .outp(out_3714)
        );        
        

        logic [WIDTH-1:0] out_3715;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.596601)
        ) inst_3715 (
            .outp(out_3715)
        );
        

        logic [WIDTH-1:0] out_3716;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3716 (
            .a(out_3715),
            .b(out_127),
            .outp(out_3716)
        );        
        

        logic [WIDTH-1:0] out_3717;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3717 (
            .a(out_3716),
            .b(out_1011),
            .outp(out_3717)
        );        
        

        logic [WIDTH-1:0] out_3718;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3718 (
            .a(out_1696),
            .b(out_3717),
            .outp(out_3718)
        );        
        

        logic [WIDTH-1:0] out_3719;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4066)
        ) inst_3719 (
            .outp(out_3719)
        );
        

        logic [WIDTH-1:0] out_3720;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3720 (
            .a(out_3719),
            .b(out_127),
            .outp(out_3720)
        );        
        

        logic [WIDTH-1:0] out_3721;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3721 (
            .a(out_1017),
            .b(out_3720),
            .outp(out_3721)
        );        
        

        logic [WIDTH-1:0] out_3722;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3722 (
            .a(out_3718),
            .b(out_3721),
            .outp(out_3722)
        );        
        

        logic [WIDTH-1:0] out_3723;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3723 (
            .a(out_3714),
            .b(out_3722),
            .outp(out_3723)
        );        
        

        logic [WIDTH-1:0] out_3724;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3724 (
            .a(out_3720),
            .b(out_1017),
            .outp(out_3724)
        );        
        

        logic [WIDTH-1:0] out_3725;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3725 (
            .a(out_1695),
            .b(out_3724),
            .outp(out_3725)
        );        
        

        logic [WIDTH-1:0] out_3726;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3726 (
            .a(out_1011),
            .b(out_3716),
            .outp(out_3726)
        );        
        

        logic [WIDTH-1:0] out_3727;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3727 (
            .a(out_3725),
            .b(out_3726),
            .outp(out_3727)
        );        
        

        logic [WIDTH-1:0] out_3728;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3728 (
            .a(out_3723),
            .b(out_3727),
            .outp(out_3728)
        );        
        

        logic [WIDTH-1:0] out_3729;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3729 (
            .a(out_1714),
            .b(out_3724),
            .outp(out_3729)
        );        
        

        logic [WIDTH-1:0] out_3730;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6516)
        ) inst_3730 (
            .outp(out_3730)
        );
        

        logic [WIDTH-1:0] out_3731;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3731 (
            .a(out_3730),
            .b(out_127),
            .outp(out_3731)
        );        
        

        logic [WIDTH-1:0] out_3732;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3732 (
            .a(out_1011),
            .b(out_3731),
            .outp(out_3732)
        );        
        

        logic [WIDTH-1:0] out_3733;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3733 (
            .a(out_3729),
            .b(out_3732),
            .outp(out_3733)
        );        
        

        logic [WIDTH-1:0] out_3734;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3734 (
            .a(out_3728),
            .b(out_3733),
            .outp(out_3734)
        );        
        

        logic [WIDTH-1:0] out_3735;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3735 (
            .a(out_1723),
            .b(out_3721),
            .outp(out_3735)
        );        
        

        logic [WIDTH-1:0] out_3736;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3736 (
            .a(out_3731),
            .b(out_1011),
            .outp(out_3736)
        );        
        

        logic [WIDTH-1:0] out_3737;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3737 (
            .a(out_3735),
            .b(out_3736),
            .outp(out_3737)
        );        
        

        logic [WIDTH-1:0] out_3738;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3738 (
            .a(out_3734),
            .b(out_3737),
            .outp(out_3738)
        );        
        

        logic [WIDTH-1:0] out_3739;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5966)
        ) inst_3739 (
            .outp(out_3739)
        );
        

        logic [WIDTH-1:0] out_3740;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3740 (
            .a(out_3739),
            .b(out_127),
            .outp(out_3740)
        );        
        

        logic [WIDTH-1:0] out_3741;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3741 (
            .a(out_3740),
            .b(out_1011),
            .outp(out_3741)
        );        
        

        logic [WIDTH-1:0] out_3742;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3742 (
            .a(out_1727),
            .b(out_3741),
            .outp(out_3742)
        );        
        

        logic [WIDTH-1:0] out_3743;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.461601)
        ) inst_3743 (
            .outp(out_3743)
        );
        

        logic [WIDTH-1:0] out_3744;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3744 (
            .a(out_3743),
            .b(out_127),
            .outp(out_3744)
        );        
        

        logic [WIDTH-1:0] out_3745;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3745 (
            .a(out_1017),
            .b(out_3744),
            .outp(out_3745)
        );        
        

        logic [WIDTH-1:0] out_3746;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3746 (
            .a(out_3742),
            .b(out_3745),
            .outp(out_3746)
        );        
        

        logic [WIDTH-1:0] out_3747;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3747 (
            .a(out_3738),
            .b(out_3746),
            .outp(out_3747)
        );        
        

        logic [WIDTH-1:0] out_3748;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3748 (
            .a(out_1726),
            .b(out_3726),
            .outp(out_3748)
        );        
        

        logic [WIDTH-1:0] out_3749;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3749 (
            .a(out_3744),
            .b(out_1017),
            .outp(out_3749)
        );        
        

        logic [WIDTH-1:0] out_3750;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3750 (
            .a(out_3748),
            .b(out_3749),
            .outp(out_3750)
        );        
        

        logic [WIDTH-1:0] out_3751;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3751 (
            .a(out_3747),
            .b(out_3750),
            .outp(out_3751)
        );        
        

        logic [WIDTH-1:0] out_3752;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3752 (
            .a(out_1740),
            .b(out_3732),
            .outp(out_3752)
        );        
        

        logic [WIDTH-1:0] out_3753;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3753 (
            .a(out_3752),
            .b(out_3749),
            .outp(out_3753)
        );        
        

        logic [WIDTH-1:0] out_3754;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3754 (
            .a(out_3751),
            .b(out_3753),
            .outp(out_3754)
        );        
        

        logic [WIDTH-1:0] out_3755;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3755 (
            .a(out_1744),
            .b(out_3736),
            .outp(out_3755)
        );        
        

        logic [WIDTH-1:0] out_3756;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3756 (
            .a(out_3755),
            .b(out_3745),
            .outp(out_3756)
        );        
        

        logic [WIDTH-1:0] out_3757;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3757 (
            .a(out_3754),
            .b(out_3756),
            .outp(out_3757)
        );        
        

        logic [WIDTH-1:0] out_3758;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5066)
        ) inst_3758 (
            .outp(out_3758)
        );
        

        logic [WIDTH-1:0] out_3759;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3759 (
            .a(out_3758),
            .b(out_1011),
            .outp(out_3759)
        );        
        

        logic [WIDTH-1:0] out_3760;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3760 (
            .a(out_3759),
            .b(out_127),
            .outp(out_3760)
        );        
        

        logic [WIDTH-1:0] out_3761;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3761 (
            .in(out_3760),
            .outp(out_3761)
        );
        

        logic [WIDTH-1:0] out_3762;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3762 (
            .a(out_1727),
            .b(out_3761),
            .outp(out_3762)
        );        
        

        logic [WIDTH-1:0] out_3763;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.6416)
        ) inst_3763 (
            .outp(out_3763)
        );
        

        logic [WIDTH-1:0] out_3764;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3764 (
            .a(out_3763),
            .b(out_1017),
            .outp(out_3764)
        );        
        

        logic [WIDTH-1:0] out_3765;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3765 (
            .a(out_3764),
            .b(out_127),
            .outp(out_3765)
        );        
        

        logic [WIDTH-1:0] out_3766;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3766 (
            .a(out_3762),
            .b(out_3765),
            .outp(out_3766)
        );        
        

        logic [WIDTH-1:0] out_3767;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3767 (
            .a(out_3757),
            .b(out_3766),
            .outp(out_3767)
        );        
        

        logic [WIDTH-1:0] out_3768;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3768 (
            .in(out_3765),
            .outp(out_3768)
        );
        

        logic [WIDTH-1:0] out_3769;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3769 (
            .a(out_1726),
            .b(out_3768),
            .outp(out_3769)
        );        
        

        logic [WIDTH-1:0] out_3770;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5066)
        ) inst_3770 (
            .outp(out_3770)
        );
        

        logic [WIDTH-1:0] out_3771;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3771 (
            .a(out_3770),
            .b(out_1011),
            .outp(out_3771)
        );        
        

        logic [WIDTH-1:0] out_3772;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3772 (
            .a(out_3771),
            .b(out_127),
            .outp(out_3772)
        );        
        

        logic [WIDTH-1:0] out_3773;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3773 (
            .a(out_3769),
            .b(out_3772),
            .outp(out_3773)
        );        
        

        logic [WIDTH-1:0] out_3774;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3774 (
            .a(out_3767),
            .b(out_3773),
            .outp(out_3774)
        );        
        

        logic [WIDTH-1:0] out_3775;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3775 (
            .a(out_1740),
            .b(out_3768),
            .outp(out_3775)
        );        
        

        logic [WIDTH-1:0] out_3776;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.4516)
        ) inst_3776 (
            .outp(out_3776)
        );
        

        logic [WIDTH-1:0] out_3777;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3777 (
            .a(out_3776),
            .b(out_1011),
            .outp(out_3777)
        );        
        

        logic [WIDTH-1:0] out_3778;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3778 (
            .a(out_3777),
            .b(out_127),
            .outp(out_3778)
        );        
        

        logic [WIDTH-1:0] out_3779;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3779 (
            .a(out_3775),
            .b(out_3778),
            .outp(out_3779)
        );        
        

        logic [WIDTH-1:0] out_3780;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3780 (
            .a(out_3774),
            .b(out_3779),
            .outp(out_3780)
        );        
        

        logic [WIDTH-1:0] out_3781;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3781 (
            .a(out_1744),
            .b(out_3765),
            .outp(out_3781)
        );        
        

        logic [WIDTH-1:0] out_3782;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3782 (
            .in(out_3778),
            .outp(out_3782)
        );
        

        logic [WIDTH-1:0] out_3783;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3783 (
            .a(out_3781),
            .b(out_3782),
            .outp(out_3783)
        );        
        

        logic [WIDTH-1:0] out_3784;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3784 (
            .a(out_3780),
            .b(out_3783),
            .outp(out_3784)
        );        
        

        logic [WIDTH-1:0] out_3785;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.3305)
        ) inst_3785 (
            .outp(out_3785)
        );
        

        logic [WIDTH-1:0] out_3786;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3786 (
            .a(out_3),
            .b(out_3785),
            .outp(out_3786)
        );        
        

        logic [WIDTH-1:0] out_3787;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3787 (
            .a(out_2072),
            .b(out_3786),
            .outp(out_3787)
        );        
        

        logic [WIDTH-1:0] out_3788;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.9305)
        ) inst_3788 (
            .outp(out_3788)
        );
        

        logic [WIDTH-1:0] out_3789;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3789 (
            .a(out_3788),
            .b(out_3),
            .outp(out_3789)
        );        
        

        logic [WIDTH-1:0] out_3790;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3790 (
            .a(out_3787),
            .b(out_3789),
            .outp(out_3790)
        );        
        

        logic [WIDTH-1:0] out_3791;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3791 (
            .a(out_3784),
            .b(out_3790),
            .outp(out_3791)
        );        
        

        logic [WIDTH-1:0] out_3792;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3792 (
            .a(out_1860),
            .b(out_1975),
            .outp(out_3792)
        );        
        

        logic [WIDTH-1:0] out_3793;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3793 (
            .a(out_3792),
            .b(out_3786),
            .outp(out_3793)
        );        
        

        logic [WIDTH-1:0] out_3794;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3794 (
            .a(out_3793),
            .b(out_3789),
            .outp(out_3794)
        );        
        

        logic [WIDTH-1:0] out_3795;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3795 (
            .in(out_3786),
            .outp(out_3795)
        );
        

        logic [WIDTH-1:0] out_3796;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3796 (
            .a(out_1977),
            .b(out_3795),
            .outp(out_3796)
        );        
        

        logic [WIDTH-1:0] out_3797;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3797 (
            .in(out_3796),
            .outp(out_3797)
        );
        

        logic [WIDTH-1:0] out_3798;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3798 (
            .a(out_336),
            .b(out_3797),
            .outp(out_3798)
        );        
        

        logic [WIDTH-1:0] out_3799;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3799 (
            .a(out_3794),
            .b(out_3798),
            .outp(out_3799)
        );        
        

        logic [WIDTH-1:0] out_3800;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3800 (
            .a(out_3797),
            .b(out_343),
            .outp(out_3800)
        );        
        

        logic [WIDTH-1:0] out_3801;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3801 (
            .a(out_3799),
            .b(out_3800),
            .outp(out_3801)
        );        
        

        logic [WIDTH-1:0] out_3802;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3802 (
            .a(out_3791),
            .b(out_3801),
            .outp(out_3802)
        );        
        

        logic [WIDTH-1:0] out_3803;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.55)
        ) inst_3803 (
            .outp(out_3803)
        );
        

        logic [WIDTH-1:0] out_3804;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3804 (
            .a(out_3803),
            .b(out_14),
            .outp(out_3804)
        );        
        

        logic [WIDTH-1:0] out_3805;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3805 (
            .a(out_1660),
            .b(out_3804),
            .outp(out_3805)
        );        
        

        logic [WIDTH-1:0] out_3806;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.8105)
        ) inst_3806 (
            .outp(out_3806)
        );
        

        logic [WIDTH-1:0] out_3807;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3807 (
            .a(out_3),
            .b(out_3806),
            .outp(out_3807)
        );        
        

        logic [WIDTH-1:0] out_3808;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3808 (
            .a(out_3805),
            .b(out_3807),
            .outp(out_3808)
        );        
        

        logic [WIDTH-1:0] out_3809;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.7105)
        ) inst_3809 (
            .outp(out_3809)
        );
        

        logic [WIDTH-1:0] out_3810;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3810 (
            .a(out_3809),
            .b(out_3),
            .outp(out_3810)
        );        
        

        logic [WIDTH-1:0] out_3811;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3811 (
            .a(out_3808),
            .b(out_3810),
            .outp(out_3811)
        );        
        

        logic [WIDTH-1:0] out_3812;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3812 (
            .a(out_3802),
            .b(out_3811),
            .outp(out_3812)
        );        
        

        logic [WIDTH-1:0] out_3813;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.993357)
        ) inst_3813 (
            .outp(out_3813)
        );
        

        logic [WIDTH-1:0] out_3814;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3814 (
            .a(out_3813),
            .b(out_1495),
            .outp(out_3814)
        );        
        

        logic [WIDTH-1:0] out_3815;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3815 (
            .a(out_3),
            .b(out_3814),
            .outp(out_3815)
        );        
        

        logic [WIDTH-1:0] out_3816;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3816 (
            .in(out_3815),
            .outp(out_3816)
        );
        

        logic [WIDTH-1:0] out_3817;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3817 (
            .a(out_1873),
            .b(out_3816),
            .outp(out_3817)
        );        
        

        logic [WIDTH-1:0] out_3818;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3818 (
            .in(out_3817),
            .outp(out_3818)
        );
        

        logic [WIDTH-1:0] out_3819;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3819 (
            .a(out_9),
            .b(out_3818),
            .outp(out_3819)
        );        
        

        logic [WIDTH-1:0] out_3820;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3820 (
            .a(out_3818),
            .b(out_21),
            .outp(out_3820)
        );        
        

        logic [WIDTH-1:0] out_3821;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3821 (
            .a(out_3819),
            .b(out_3820),
            .outp(out_3821)
        );        
        

        logic [WIDTH-1:0] out_3822;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3822 (
            .a(out_3812),
            .b(out_3821),
            .outp(out_3822)
        );        
        

        logic [WIDTH-1:0] out_3823;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.000499725)
        ) inst_3823 (
            .outp(out_3823)
        );
        

        logic [WIDTH-1:0] out_3824;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3824 (
            .a(out_3),
            .b(out_3823),
            .outp(out_3824)
        );        
        

        logic [WIDTH-1:0] out_3825;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3825 (
            .a(out_1862),
            .b(out_3824),
            .outp(out_3825)
        );        
        

        logic [WIDTH-1:0] out_3826;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0995007)
        ) inst_3826 (
            .outp(out_3826)
        );
        

        logic [WIDTH-1:0] out_3827;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3827 (
            .a(out_3826),
            .b(out_3),
            .outp(out_3827)
        );        
        

        logic [WIDTH-1:0] out_3828;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3828 (
            .in(out_3827),
            .outp(out_3828)
        );
        

        logic [WIDTH-1:0] out_3829;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3829 (
            .a(out_3825),
            .b(out_3828),
            .outp(out_3829)
        );        
        

        logic [WIDTH-1:0] out_3830;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3830 (
            .a(out_3822),
            .b(out_3829),
            .outp(out_3830)
        );        
        

        logic [WIDTH-1:0] out_3831;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.150499)
        ) inst_3831 (
            .outp(out_3831)
        );
        

        logic [WIDTH-1:0] out_3832;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3832 (
            .a(out_3),
            .b(out_3831),
            .outp(out_3832)
        );        
        

        logic [WIDTH-1:0] out_3833;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3833 (
            .a(out_1649),
            .b(out_3832),
            .outp(out_3833)
        );        
        

        logic [WIDTH-1:0] out_3834;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.249501)
        ) inst_3834 (
            .outp(out_3834)
        );
        

        logic [WIDTH-1:0] out_3835;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3835 (
            .a(out_3834),
            .b(out_3),
            .outp(out_3835)
        );        
        

        logic [WIDTH-1:0] out_3836;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3836 (
            .in(out_3835),
            .outp(out_3836)
        );
        

        logic [WIDTH-1:0] out_3837;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3837 (
            .a(out_3833),
            .b(out_3836),
            .outp(out_3837)
        );        
        

        logic [WIDTH-1:0] out_3838;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3838 (
            .a(out_3830),
            .b(out_3837),
            .outp(out_3838)
        );        
        

        logic [WIDTH-1:0] out_3839;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3839 (
            .a(out_1660),
            .b(out_1663),
            .outp(out_3839)
        );        
        

        logic [WIDTH-1:0] out_3840;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3840 (
            .a(out_3839),
            .b(out_3832),
            .outp(out_3840)
        );        
        

        logic [WIDTH-1:0] out_3841;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3841 (
            .a(out_3840),
            .b(out_3836),
            .outp(out_3841)
        );        
        

        logic [WIDTH-1:0] out_3842;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3842 (
            .in(out_3832),
            .outp(out_3842)
        );
        

        logic [WIDTH-1:0] out_3843;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3843 (
            .a(out_1664),
            .b(out_3842),
            .outp(out_3843)
        );        
        

        logic [WIDTH-1:0] out_3844;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3844 (
            .in(out_3843),
            .outp(out_3844)
        );
        

        logic [WIDTH-1:0] out_3845;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3845 (
            .a(out_336),
            .b(out_3844),
            .outp(out_3845)
        );        
        

        logic [WIDTH-1:0] out_3846;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3846 (
            .a(out_3841),
            .b(out_3845),
            .outp(out_3846)
        );        
        

        logic [WIDTH-1:0] out_3847;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3847 (
            .a(out_3844),
            .b(out_343),
            .outp(out_3847)
        );        
        

        logic [WIDTH-1:0] out_3848;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3848 (
            .a(out_3846),
            .b(out_3847),
            .outp(out_3848)
        );        
        

        logic [WIDTH-1:0] out_3849;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3849 (
            .a(out_3838),
            .b(out_3848),
            .outp(out_3849)
        );        
        

        logic [WIDTH-1:0] out_3850;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.66785)
        ) inst_3850 (
            .outp(out_3850)
        );
        

        logic [WIDTH-1:0] out_3851;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3851 (
            .a(out_3850),
            .b(out_127),
            .outp(out_3851)
        );        
        

        logic [WIDTH-1:0] out_3852;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3852 (
            .a(out_3851),
            .b(out_928),
            .outp(out_3852)
        );        
        

        logic [WIDTH-1:0] out_3853;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.24785)
        ) inst_3853 (
            .outp(out_3853)
        );
        

        logic [WIDTH-1:0] out_3854;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3854 (
            .a(out_3853),
            .b(out_127),
            .outp(out_3854)
        );        
        

        logic [WIDTH-1:0] out_3855;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3855 (
            .in(out_3854),
            .outp(out_3855)
        );
        

        logic [WIDTH-1:0] out_3856;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3856 (
            .a(out_3852),
            .b(out_3855),
            .outp(out_3856)
        );        
        

        logic [WIDTH-1:0] out_3857;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.36)
        ) inst_3857 (
            .outp(out_3857)
        );
        

        logic [WIDTH-1:0] out_3858;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3858 (
            .a(out_3857),
            .b(out_928),
            .outp(out_3858)
        );        
        

        logic [WIDTH-1:0] out_3859;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3859 (
            .a(out_3856),
            .b(out_3858),
            .outp(out_3859)
        );        
        

        logic [WIDTH-1:0] out_3860;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3860 (
            .a(out_928),
            .b(out_3851),
            .outp(out_3860)
        );        
        

        logic [WIDTH-1:0] out_3861;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3861 (
            .a(out_3854),
            .b(out_3860),
            .outp(out_3861)
        );        
        

        logic [WIDTH-1:0] out_3862;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3862 (
            .in(out_3858),
            .outp(out_3862)
        );
        

        logic [WIDTH-1:0] out_3863;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3863 (
            .a(out_3861),
            .b(out_3862),
            .outp(out_3863)
        );        
        

        logic [WIDTH-1:0] out_3864;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3864 (
            .a(out_3859),
            .b(out_3863),
            .outp(out_3864)
        );        
        

        logic [WIDTH-1:0] out_3865;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3865 (
            .a(out_2943),
            .b(out_566),
            .outp(out_3865)
        );        
        

        logic [WIDTH-1:0] out_3866;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.7935)
        ) inst_3866 (
            .outp(out_3866)
        );
        

        logic [WIDTH-1:0] out_3867;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3867 (
            .a(out_3866),
            .b(out_862),
            .outp(out_3867)
        );        
        

        logic [WIDTH-1:0] out_3868;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3868 (
            .a(out_3865),
            .b(out_3867),
            .outp(out_3868)
        );        
        

        logic [WIDTH-1:0] out_3869;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.4935)
        ) inst_3869 (
            .outp(out_3869)
        );
        

        logic [WIDTH-1:0] out_3870;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3870 (
            .a(out_3869),
            .b(out_868),
            .outp(out_3870)
        );        
        

        logic [WIDTH-1:0] out_3871;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3871 (
            .in(out_3870),
            .outp(out_3871)
        );
        

        logic [WIDTH-1:0] out_3872;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3872 (
            .a(out_3868),
            .b(out_3871),
            .outp(out_3872)
        );        
        

        logic [WIDTH-1:0] out_3873;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3873 (
            .a(out_3864),
            .b(out_3872),
            .outp(out_3873)
        );        
        

        logic [WIDTH-1:0] out_3874;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3874 (
            .in(out_3867),
            .outp(out_3874)
        );
        

        logic [WIDTH-1:0] out_3875;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3875 (
            .a(out_3870),
            .b(out_3874),
            .outp(out_3875)
        );        
        

        logic [WIDTH-1:0] out_3876;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3876 (
            .in(out_3865),
            .outp(out_3876)
        );
        

        logic [WIDTH-1:0] out_3877;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3877 (
            .a(out_3875),
            .b(out_3876),
            .outp(out_3877)
        );        
        

        logic [WIDTH-1:0] out_3878;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3878 (
            .a(out_3873),
            .b(out_3877),
            .outp(out_3878)
        );        
        

        logic [WIDTH-1:0] out_3879;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.497)
        ) inst_3879 (
            .outp(out_3879)
        );
        

        logic [WIDTH-1:0] out_3880;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3880 (
            .a(out_3879),
            .b(out_3),
            .outp(out_3880)
        );        
        

        logic [WIDTH-1:0] out_3881;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3881 (
            .a(out_3880),
            .b(out_878),
            .outp(out_3881)
        );        
        

        logic [WIDTH-1:0] out_3882;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.89845)
        ) inst_3882 (
            .outp(out_3882)
        );
        

        logic [WIDTH-1:0] out_3883;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3883 (
            .a(out_3882),
            .b(out_884),
            .outp(out_3883)
        );        
        

        logic [WIDTH-1:0] out_3884;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3884 (
            .a(out_3883),
            .b(out_886),
            .outp(out_3884)
        );        
        

        logic [WIDTH-1:0] out_3885;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3885 (
            .in(out_3884),
            .outp(out_3885)
        );
        

        logic [WIDTH-1:0] out_3886;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3886 (
            .a(out_3881),
            .b(out_3885),
            .outp(out_3886)
        );        
        

        logic [WIDTH-1:0] out_3887;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.95355)
        ) inst_3887 (
            .outp(out_3887)
        );
        

        logic [WIDTH-1:0] out_3888;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3888 (
            .a(out_3887),
            .b(out_894),
            .outp(out_3888)
        );        
        

        logic [WIDTH-1:0] out_3889;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3889 (
            .a(out_891),
            .b(out_3888),
            .outp(out_3889)
        );        
        

        logic [WIDTH-1:0] out_3890;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3890 (
            .a(out_3886),
            .b(out_3889),
            .outp(out_3890)
        );        
        

        logic [WIDTH-1:0] out_3891;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3891 (
            .a(out_3878),
            .b(out_3890),
            .outp(out_3891)
        );        
        

        logic [WIDTH-1:0] out_3892;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3892 (
            .a(out_3888),
            .b(out_891),
            .outp(out_3892)
        );        
        

        logic [WIDTH-1:0] out_3893;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.89845)
        ) inst_3893 (
            .outp(out_3893)
        );
        

        logic [WIDTH-1:0] out_3894;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3894 (
            .a(out_3893),
            .b(out_884),
            .outp(out_3894)
        );        
        

        logic [WIDTH-1:0] out_3895;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3895 (
            .a(out_3894),
            .b(out_886),
            .outp(out_3895)
        );        
        

        logic [WIDTH-1:0] out_3896;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3896 (
            .a(out_3892),
            .b(out_3895),
            .outp(out_3896)
        );        
        

        logic [WIDTH-1:0] out_3897;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3897 (
            .a(out_878),
            .b(out_3880),
            .outp(out_3897)
        );        
        

        logic [WIDTH-1:0] out_3898;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3898 (
            .a(out_3896),
            .b(out_3897),
            .outp(out_3898)
        );        
        

        logic [WIDTH-1:0] out_3899;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3899 (
            .a(out_3891),
            .b(out_3898),
            .outp(out_3899)
        );        
        

        logic [WIDTH-1:0] out_3900;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.54)
        ) inst_3900 (
            .outp(out_3900)
        );
        

        logic [WIDTH-1:0] out_3901;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3901 (
            .a(out_3900),
            .b(out_910),
            .outp(out_3901)
        );        
        

        logic [WIDTH-1:0] out_3902;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3902 (
            .in(out_3901),
            .outp(out_3902)
        );
        

        logic [WIDTH-1:0] out_3903;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.43045)
        ) inst_3903 (
            .outp(out_3903)
        );
        

        logic [WIDTH-1:0] out_3904;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3904 (
            .a(out_3903),
            .b(out_886),
            .outp(out_3904)
        );        
        

        logic [WIDTH-1:0] out_3905;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3905 (
            .in(out_3904),
            .outp(out_3905)
        );
        

        logic [WIDTH-1:0] out_3906;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3906 (
            .a(out_3902),
            .b(out_3905),
            .outp(out_3906)
        );        
        

        logic [WIDTH-1:0] out_3907;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.87595)
        ) inst_3907 (
            .outp(out_3907)
        );
        

        logic [WIDTH-1:0] out_3908;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3908 (
            .a(out_3907),
            .b(out_910),
            .outp(out_3908)
        );        
        

        logic [WIDTH-1:0] out_3909;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3909 (
            .a(out_3908),
            .b(out_886),
            .outp(out_3909)
        );        
        

        logic [WIDTH-1:0] out_3910;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3910 (
            .a(out_3906),
            .b(out_3909),
            .outp(out_3910)
        );        
        

        logic [WIDTH-1:0] out_3911;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3911 (
            .a(out_3899),
            .b(out_3910),
            .outp(out_3911)
        );        
        

        logic [WIDTH-1:0] out_3912;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3912 (
            .a(out_3901),
            .b(out_3904),
            .outp(out_3912)
        );        
        

        logic [WIDTH-1:0] out_3913;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3913 (
            .in(out_3909),
            .outp(out_3913)
        );
        

        logic [WIDTH-1:0] out_3914;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3914 (
            .a(out_3912),
            .b(out_3913),
            .outp(out_3914)
        );        
        

        logic [WIDTH-1:0] out_3915;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3915 (
            .a(out_3911),
            .b(out_3914),
            .outp(out_3915)
        );        
        

        logic [WIDTH-1:0] out_3916;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3916 (
            .in(out_3915),
            .outp(out_3916)
        );
        

        logic [WIDTH-1:0] out_3917;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3917 (
            .a(out_1870),
            .b(out_3916),
            .outp(out_3917)
        );        
        

        logic [WIDTH-1:0] out_3918;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.687)
        ) inst_3918 (
            .outp(out_3918)
        );
        

        logic [WIDTH-1:0] out_3919;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3919 (
            .a(out_3918),
            .b(out_3),
            .outp(out_3919)
        );        
        

        logic [WIDTH-1:0] out_3920;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3920 (
            .a(out_3917),
            .b(out_3919),
            .outp(out_3920)
        );        
        

        logic [WIDTH-1:0] out_3921;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.187)
        ) inst_3921 (
            .outp(out_3921)
        );
        

        logic [WIDTH-1:0] out_3922;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3922 (
            .a(out_3921),
            .b(out_3),
            .outp(out_3922)
        );        
        

        logic [WIDTH-1:0] out_3923;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3923 (
            .in(out_3922),
            .outp(out_3923)
        );
        

        logic [WIDTH-1:0] out_3924;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3924 (
            .a(out_3920),
            .b(out_3923),
            .outp(out_3924)
        );        
        

        logic [WIDTH-1:0] out_3925;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3925 (
            .a(out_3849),
            .b(out_3924),
            .outp(out_3925)
        );        
        

        logic [WIDTH-1:0] out_3926;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.307)
        ) inst_3926 (
            .outp(out_3926)
        );
        

        logic [WIDTH-1:0] out_3927;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3927 (
            .a(out_3926),
            .b(out_3),
            .outp(out_3927)
        );        
        

        logic [WIDTH-1:0] out_3928;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3928 (
            .a(out_3805),
            .b(out_3927),
            .outp(out_3928)
        );        
        

        logic [WIDTH-1:0] out_3929;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.407)
        ) inst_3929 (
            .outp(out_3929)
        );
        

        logic [WIDTH-1:0] out_3930;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3930 (
            .a(out_3929),
            .b(out_3),
            .outp(out_3930)
        );        
        

        logic [WIDTH-1:0] out_3931;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3931 (
            .in(out_3930),
            .outp(out_3931)
        );
        

        logic [WIDTH-1:0] out_3932;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3932 (
            .a(out_3928),
            .b(out_3931),
            .outp(out_3932)
        );        
        

        logic [WIDTH-1:0] out_3933;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3933 (
            .a(out_3925),
            .b(out_3932),
            .outp(out_3933)
        );        
        

        logic [WIDTH-1:0] out_3934;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.12414)
        ) inst_3934 (
            .outp(out_3934)
        );
        

        logic [WIDTH-1:0] out_3935;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3935 (
            .a(out_3934),
            .b(out_3),
            .outp(out_3935)
        );        
        

        logic [WIDTH-1:0] out_3936;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3936 (
            .a(out_3935),
            .b(out_1495),
            .outp(out_3936)
        );        
        

        logic [WIDTH-1:0] out_3937;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3937 (
            .in(out_3936),
            .outp(out_3937)
        );
        

        logic [WIDTH-1:0] out_3938;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3938 (
            .a(out_1873),
            .b(out_3937),
            .outp(out_3938)
        );        
        

        logic [WIDTH-1:0] out_3939;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3939 (
            .in(out_3938),
            .outp(out_3939)
        );
        

        logic [WIDTH-1:0] out_3940;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3940 (
            .a(out_9),
            .b(out_3939),
            .outp(out_3940)
        );        
        

        logic [WIDTH-1:0] out_3941;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3941 (
            .a(out_3939),
            .b(out_21),
            .outp(out_3941)
        );        
        

        logic [WIDTH-1:0] out_3942;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3942 (
            .a(out_3940),
            .b(out_3941),
            .outp(out_3942)
        );        
        

        logic [WIDTH-1:0] out_3943;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3943 (
            .a(out_3933),
            .b(out_3942),
            .outp(out_3943)
        );        
        

        logic [WIDTH-1:0] out_3944;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.585)
        ) inst_3944 (
            .outp(out_3944)
        );
        

        logic [WIDTH-1:0] out_3945;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3945 (
            .a(out_3944),
            .b(out_14),
            .outp(out_3945)
        );        
        

        logic [WIDTH-1:0] out_3946;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.675)
        ) inst_3946 (
            .outp(out_3946)
        );
        

        logic [WIDTH-1:0] out_3947;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3947 (
            .a(out_3946),
            .b(out_14),
            .outp(out_3947)
        );        
        

        logic [WIDTH-1:0] out_3948;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3948 (
            .in(out_3947),
            .outp(out_3948)
        );
        

        logic [WIDTH-1:0] out_3949;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3949 (
            .a(out_3945),
            .b(out_3948),
            .outp(out_3949)
        );        
        

        logic [WIDTH-1:0] out_3950;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.967)
        ) inst_3950 (
            .outp(out_3950)
        );
        

        logic [WIDTH-1:0] out_3951;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3951 (
            .a(out_3950),
            .b(out_3),
            .outp(out_3951)
        );        
        

        logic [WIDTH-1:0] out_3952;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3952 (
            .a(out_3949),
            .b(out_3951),
            .outp(out_3952)
        );        
        

        logic [WIDTH-1:0] out_3953;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.467)
        ) inst_3953 (
            .outp(out_3953)
        );
        

        logic [WIDTH-1:0] out_3954;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3954 (
            .a(out_3953),
            .b(out_3),
            .outp(out_3954)
        );        
        

        logic [WIDTH-1:0] out_3955;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3955 (
            .in(out_3954),
            .outp(out_3955)
        );
        

        logic [WIDTH-1:0] out_3956;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3956 (
            .a(out_3952),
            .b(out_3955),
            .outp(out_3956)
        );        
        

        logic [WIDTH-1:0] out_3957;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.242)
        ) inst_3957 (
            .outp(out_3957)
        );
        

        logic [WIDTH-1:0] out_3958;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3958 (
            .a(out_3957),
            .b(out_3),
            .outp(out_3958)
        );        
        

        logic [WIDTH-1:0] out_3959;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3959 (
            .in(out_3958),
            .outp(out_3959)
        );
        

        logic [WIDTH-1:0] out_3960;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3960 (
            .a(out_1873),
            .b(out_3959),
            .outp(out_3960)
        );        
        

        logic [WIDTH-1:0] out_3961;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3961 (
            .in(out_3960),
            .outp(out_3961)
        );
        

        logic [WIDTH-1:0] out_3962;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3962 (
            .a(out_3961),
            .b(out_21),
            .outp(out_3962)
        );        
        

        logic [WIDTH-1:0] out_3963;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.05625)
        ) inst_3963 (
            .outp(out_3963)
        );
        

        logic [WIDTH-1:0] out_3964;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3964 (
            .a(out_3963),
            .b(out_553),
            .outp(out_3964)
        );        
        

        logic [WIDTH-1:0] out_3965;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.06718)
        ) inst_3965 (
            .outp(out_3965)
        );
        

        logic [WIDTH-1:0] out_3966;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3966 (
            .a(out_3965),
            .b(out_556),
            .outp(out_3966)
        );        
        

        logic [WIDTH-1:0] out_3967;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3967 (
            .a(out_3966),
            .b(out_559),
            .outp(out_3967)
        );        
        

        logic [WIDTH-1:0] out_3968;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3968 (
            .a(out_3964),
            .b(out_3967),
            .outp(out_3968)
        );        
        

        logic [WIDTH-1:0] out_3969;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.30217)
        ) inst_3969 (
            .outp(out_3969)
        );
        

        logic [WIDTH-1:0] out_3970;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3970 (
            .a(out_556),
            .b(out_3969),
            .outp(out_3970)
        );        
        

        logic [WIDTH-1:0] out_3971;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3971 (
            .a(out_3970),
            .b(out_566),
            .outp(out_3971)
        );        
        

        logic [WIDTH-1:0] out_3972;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3972 (
            .in(out_3971),
            .outp(out_3972)
        );
        

        logic [WIDTH-1:0] out_3973;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3973 (
            .a(out_3968),
            .b(out_3972),
            .outp(out_3973)
        );        
        

        logic [WIDTH-1:0] out_3974;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3974 (
            .a(out_559),
            .b(out_3966),
            .outp(out_3974)
        );        
        

        logic [WIDTH-1:0] out_3975;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3975 (
            .a(out_3971),
            .b(out_3974),
            .outp(out_3975)
        );        
        

        logic [WIDTH-1:0] out_3976;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3976 (
            .in(out_3964),
            .outp(out_3976)
        );
        

        logic [WIDTH-1:0] out_3977;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3977 (
            .a(out_3975),
            .b(out_3976),
            .outp(out_3977)
        );        
        

        logic [WIDTH-1:0] out_3978;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3978 (
            .a(out_3973),
            .b(out_3977),
            .outp(out_3978)
        );        
        

        logic [WIDTH-1:0] out_3979;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3979 (
            .in(out_3978),
            .outp(out_3979)
        );
        

        logic [WIDTH-1:0] out_3980;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3980 (
            .a(out_3962),
            .b(out_3979),
            .outp(out_3980)
        );        
        

        logic [WIDTH-1:0] out_3981;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3981 (
            .a(out_9),
            .b(out_3961),
            .outp(out_3981)
        );        
        

        logic [WIDTH-1:0] out_3982;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3982 (
            .a(out_3980),
            .b(out_3981),
            .outp(out_3982)
        );        
        

        logic [WIDTH-1:0] out_3983;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3983 (
            .a(out_3956),
            .b(out_3982),
            .outp(out_3983)
        );        
        

        logic [WIDTH-1:0] out_3984;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3984 (
            .a(out_3962),
            .b(out_3983),
            .outp(out_3984)
        );        
        

        logic [WIDTH-1:0] out_3985;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3985 (
            .a(out_3943),
            .b(out_3984),
            .outp(out_3985)
        );        
        

        logic [WIDTH-1:0] out_3986;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.875)
        ) inst_3986 (
            .outp(out_3986)
        );
        

        logic [WIDTH-1:0] out_3987;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3987 (
            .a(out_3986),
            .b(out_3),
            .outp(out_3987)
        );        
        

        logic [WIDTH-1:0] out_3988;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3988 (
            .a(out_1676),
            .b(out_3987),
            .outp(out_3988)
        );        
        

        logic [WIDTH-1:0] out_3989;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3989 (
            .in(out_3241),
            .outp(out_3989)
        );
        

        logic [WIDTH-1:0] out_3990;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3990 (
            .a(out_3988),
            .b(out_3989),
            .outp(out_3990)
        );        
        

        logic [WIDTH-1:0] out_3991;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3991 (
            .a(out_3985),
            .b(out_3990),
            .outp(out_3991)
        );        
        

        logic [WIDTH-1:0] out_3992;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.287)
        ) inst_3992 (
            .outp(out_3992)
        );
        

        logic [WIDTH-1:0] out_3993;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3993 (
            .a(out_3992),
            .b(out_3),
            .outp(out_3993)
        );        
        

        logic [WIDTH-1:0] out_3994;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3994 (
            .a(out_1660),
            .b(out_3993),
            .outp(out_3994)
        );        
        

        logic [WIDTH-1:0] out_3995;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.387)
        ) inst_3995 (
            .outp(out_3995)
        );
        

        logic [WIDTH-1:0] out_3996;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3996 (
            .a(out_3995),
            .b(out_3),
            .outp(out_3996)
        );        
        

        logic [WIDTH-1:0] out_3997;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3997 (
            .in(out_3996),
            .outp(out_3997)
        );
        

        logic [WIDTH-1:0] out_3998;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3998 (
            .a(out_3994),
            .b(out_3997),
            .outp(out_3998)
        );        
        

        logic [WIDTH-1:0] out_3999;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_3999 (
            .a(out_3998),
            .b(out_3804),
            .outp(out_3999)
        );        
        

        logic [WIDTH-1:0] out_4000;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4000 (
            .a(out_3991),
            .b(out_3999),
            .outp(out_4000)
        );        
        

        logic [WIDTH-1:0] out_4001;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.537)
        ) inst_4001 (
            .outp(out_4001)
        );
        

        logic [WIDTH-1:0] out_4002;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4002 (
            .a(out_4001),
            .b(out_3),
            .outp(out_4002)
        );        
        

        logic [WIDTH-1:0] out_4003;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4003 (
            .a(out_3805),
            .b(out_4002),
            .outp(out_4003)
        );        
        

        logic [WIDTH-1:0] out_4004;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.637)
        ) inst_4004 (
            .outp(out_4004)
        );
        

        logic [WIDTH-1:0] out_4005;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4005 (
            .a(out_4004),
            .b(out_3),
            .outp(out_4005)
        );        
        

        logic [WIDTH-1:0] out_4006;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4006 (
            .in(out_4005),
            .outp(out_4006)
        );
        

        logic [WIDTH-1:0] out_4007;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4007 (
            .a(out_4003),
            .b(out_4006),
            .outp(out_4007)
        );        
        

        logic [WIDTH-1:0] out_4008;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4008 (
            .a(out_4000),
            .b(out_4007),
            .outp(out_4008)
        );        
        

        logic [WIDTH-1:0] out_4009;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.375)
        ) inst_4009 (
            .outp(out_4009)
        );
        

        logic [WIDTH-1:0] out_4010;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4010 (
            .a(out_4009),
            .b(out_14),
            .outp(out_4010)
        );        
        

        logic [WIDTH-1:0] out_4011;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4011 (
            .a(out_1660),
            .b(out_4010),
            .outp(out_4011)
        );        
        

        logic [WIDTH-1:0] out_4012;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.787)
        ) inst_4012 (
            .outp(out_4012)
        );
        

        logic [WIDTH-1:0] out_4013;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4013 (
            .a(out_4012),
            .b(out_3),
            .outp(out_4013)
        );        
        

        logic [WIDTH-1:0] out_4014;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4014 (
            .a(out_4011),
            .b(out_4013),
            .outp(out_4014)
        );        
        

        logic [WIDTH-1:0] out_4015;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.887)
        ) inst_4015 (
            .outp(out_4015)
        );
        

        logic [WIDTH-1:0] out_4016;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4016 (
            .a(out_4015),
            .b(out_3),
            .outp(out_4016)
        );        
        

        logic [WIDTH-1:0] out_4017;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4017 (
            .in(out_4016),
            .outp(out_4017)
        );
        

        logic [WIDTH-1:0] out_4018;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4018 (
            .a(out_4014),
            .b(out_4017),
            .outp(out_4018)
        );        
        

        logic [WIDTH-1:0] out_4019;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4019 (
            .a(out_4008),
            .b(out_4018),
            .outp(out_4019)
        );        
        

        logic [WIDTH-1:0] out_4020;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4020 (
            .a(out_1645),
            .b(out_4017),
            .outp(out_4020)
        );        
        

        logic [WIDTH-1:0] out_4021;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.55)
        ) inst_4021 (
            .outp(out_4021)
        );
        

        logic [WIDTH-1:0] out_4022;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4022 (
            .a(out_4021),
            .b(out_14),
            .outp(out_4022)
        );        
        

        logic [WIDTH-1:0] out_4023;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4023 (
            .in(out_4022),
            .outp(out_4023)
        );
        

        logic [WIDTH-1:0] out_4024;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4024 (
            .a(out_4020),
            .b(out_4023),
            .outp(out_4024)
        );        
        

        logic [WIDTH-1:0] out_4025;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.237)
        ) inst_4025 (
            .outp(out_4025)
        );
        

        logic [WIDTH-1:0] out_4026;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4026 (
            .a(out_4025),
            .b(out_3),
            .outp(out_4026)
        );        
        

        logic [WIDTH-1:0] out_4027;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4027 (
            .a(out_4024),
            .b(out_4026),
            .outp(out_4027)
        );        
        

        logic [WIDTH-1:0] out_4028;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4028 (
            .in(out_3804),
            .outp(out_4028)
        );
        

        logic [WIDTH-1:0] out_4029;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.462)
        ) inst_4029 (
            .outp(out_4029)
        );
        

        logic [WIDTH-1:0] out_4030;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4030 (
            .a(out_4029),
            .b(out_3),
            .outp(out_4030)
        );        
        

        logic [WIDTH-1:0] out_4031;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4031 (
            .in(out_4030),
            .outp(out_4031)
        );
        

        logic [WIDTH-1:0] out_4032;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4032 (
            .a(out_4028),
            .b(out_4031),
            .outp(out_4032)
        );        
        

        logic [WIDTH-1:0] out_4033;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4033 (
            .in(out_4032),
            .outp(out_4033)
        );
        

        logic [WIDTH-1:0] out_4034;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4034 (
            .a(out_460),
            .b(out_4033),
            .outp(out_4034)
        );        
        

        logic [WIDTH-1:0] out_4035;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4035 (
            .a(out_4033),
            .b(out_9),
            .outp(out_4035)
        );        
        

        logic [WIDTH-1:0] out_4036;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4036 (
            .a(out_4034),
            .b(out_4035),
            .outp(out_4036)
        );        
        

        logic [WIDTH-1:0] out_4037;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.712)
        ) inst_4037 (
            .outp(out_4037)
        );
        

        logic [WIDTH-1:0] out_4038;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4038 (
            .a(out_4037),
            .b(out_3),
            .outp(out_4038)
        );        
        

        logic [WIDTH-1:0] out_4039;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4039 (
            .in(out_4038),
            .outp(out_4039)
        );
        

        logic [WIDTH-1:0] out_4040;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4040 (
            .a(out_4028),
            .b(out_4039),
            .outp(out_4040)
        );        
        

        logic [WIDTH-1:0] out_4041;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4041 (
            .in(out_4040),
            .outp(out_4041)
        );
        

        logic [WIDTH-1:0] out_4042;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4042 (
            .a(out_460),
            .b(out_4041),
            .outp(out_4042)
        );        
        

        logic [WIDTH-1:0] out_4043;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4043 (
            .a(out_4041),
            .b(out_9),
            .outp(out_4043)
        );        
        

        logic [WIDTH-1:0] out_4044;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4044 (
            .a(out_4042),
            .b(out_4043),
            .outp(out_4044)
        );        
        

        logic [WIDTH-1:0] out_4045;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4045 (
            .a(out_4036),
            .b(out_4044),
            .outp(out_4045)
        );        
        

        logic [WIDTH-1:0] out_4046;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4046 (
            .a(out_4027),
            .b(out_4045),
            .outp(out_4046)
        );        
        

        logic [WIDTH-1:0] out_4047;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4047 (
            .a(out_4019),
            .b(out_4046),
            .outp(out_4047)
        );        
        

        logic [WIDTH-1:0] out_4048;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.89365)
        ) inst_4048 (
            .outp(out_4048)
        );
        

        logic [WIDTH-1:0] out_4049;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4049 (
            .a(out_137),
            .b(out_4048),
            .outp(out_4049)
        );        
        

        logic [WIDTH-1:0] out_4050;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4050 (
            .a(out_1891),
            .b(out_4049),
            .outp(out_4050)
        );        
        

        logic [WIDTH-1:0] out_4051;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.681276)
        ) inst_4051 (
            .outp(out_4051)
        );
        

        logic [WIDTH-1:0] out_4052;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4052 (
            .a(out_1897),
            .b(out_566),
            .outp(out_4052)
        );        
        

        logic [WIDTH-1:0] out_4053;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4053 (
            .a(out_4051),
            .b(out_4052),
            .outp(out_4053)
        );        
        

        logic [WIDTH-1:0] out_4054;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4054 (
            .a(out_4050),
            .b(out_4053),
            .outp(out_4054)
        );        
        

        logic [WIDTH-1:0] out_4055;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.01488)
        ) inst_4055 (
            .outp(out_4055)
        );
        

        logic [WIDTH-1:0] out_4056;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4056 (
            .a(out_4055),
            .b(out_1904),
            .outp(out_4056)
        );        
        

        logic [WIDTH-1:0] out_4057;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4057 (
            .a(out_4056),
            .b(out_1907),
            .outp(out_4057)
        );        
        

        logic [WIDTH-1:0] out_4058;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4058 (
            .a(out_4054),
            .b(out_4057),
            .outp(out_4058)
        );        
        

        logic [WIDTH-1:0] out_4059;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.01488)
        ) inst_4059 (
            .outp(out_4059)
        );
        

        logic [WIDTH-1:0] out_4060;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4060 (
            .a(out_4059),
            .b(out_1904),
            .outp(out_4060)
        );        
        

        logic [WIDTH-1:0] out_4061;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4061 (
            .a(out_1907),
            .b(out_4060),
            .outp(out_4061)
        );        
        

        logic [WIDTH-1:0] out_4062;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4062 (
            .a(out_4052),
            .b(out_4051),
            .outp(out_4062)
        );        
        

        logic [WIDTH-1:0] out_4063;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4063 (
            .a(out_4061),
            .b(out_4062),
            .outp(out_4063)
        );        
        

        logic [WIDTH-1:0] out_4064;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4064 (
            .a(out_4049),
            .b(out_1891),
            .outp(out_4064)
        );        
        

        logic [WIDTH-1:0] out_4065;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4065 (
            .a(out_4063),
            .b(out_4064),
            .outp(out_4065)
        );        
        

        logic [WIDTH-1:0] out_4066;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4066 (
            .a(out_4058),
            .b(out_4065),
            .outp(out_4066)
        );        
        

        logic [WIDTH-1:0] out_4067;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4067 (
            .in(out_4066),
            .outp(out_4067)
        );
        

        logic [WIDTH-1:0] out_4068;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.725)
        ) inst_4068 (
            .outp(out_4068)
        );
        

        logic [WIDTH-1:0] out_4069;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4069 (
            .a(out_4068),
            .b(out_14),
            .outp(out_4069)
        );        
        

        logic [WIDTH-1:0] out_4070;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4070 (
            .a(out_4067),
            .b(out_4069),
            .outp(out_4070)
        );        
        

        logic [WIDTH-1:0] out_4071;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.95)
        ) inst_4071 (
            .outp(out_4071)
        );
        

        logic [WIDTH-1:0] out_4072;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4072 (
            .a(out_4071),
            .b(out_14),
            .outp(out_4072)
        );        
        

        logic [WIDTH-1:0] out_4073;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4073 (
            .in(out_4072),
            .outp(out_4073)
        );
        

        logic [WIDTH-1:0] out_4074;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4074 (
            .a(out_4070),
            .b(out_4073),
            .outp(out_4074)
        );        
        

        logic [WIDTH-1:0] out_4075;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.289)
        ) inst_4075 (
            .outp(out_4075)
        );
        

        logic [WIDTH-1:0] out_4076;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4076 (
            .a(out_3),
            .b(out_4075),
            .outp(out_4076)
        );        
        

        logic [WIDTH-1:0] out_4077;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4077 (
            .a(out_4074),
            .b(out_4076),
            .outp(out_4077)
        );        
        

        logic [WIDTH-1:0] out_4078;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.139)
        ) inst_4078 (
            .outp(out_4078)
        );
        

        logic [WIDTH-1:0] out_4079;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4079 (
            .a(out_4078),
            .b(out_3),
            .outp(out_4079)
        );        
        

        logic [WIDTH-1:0] out_4080;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4080 (
            .a(out_4077),
            .b(out_4079),
            .outp(out_4080)
        );        
        

        logic [WIDTH-1:0] out_4081;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.241667)
        ) inst_4081 (
            .outp(out_4081)
        );
        

        logic [WIDTH-1:0] out_4082;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4082 (
            .a(out_4081),
            .b(out_1933),
            .outp(out_4082)
        );        
        

        logic [WIDTH-1:0] out_4083;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4083 (
            .in(out_4082),
            .outp(out_4083)
        );
        

        logic [WIDTH-1:0] out_4084;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.214)
        ) inst_4084 (
            .outp(out_4084)
        );
        

        logic [WIDTH-1:0] out_4085;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4085 (
            .a(out_3),
            .b(out_4084),
            .outp(out_4085)
        );        
        

        logic [WIDTH-1:0] out_4086;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4086 (
            .in(out_4085),
            .outp(out_4086)
        );
        

        logic [WIDTH-1:0] out_4087;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4087 (
            .a(out_4083),
            .b(out_4086),
            .outp(out_4087)
        );        
        

        logic [WIDTH-1:0] out_4088;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4088 (
            .in(out_4087),
            .outp(out_4088)
        );
        

        logic [WIDTH-1:0] out_4089;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4089 (
            .a(out_4088),
            .b(out_460),
            .outp(out_4089)
        );        
        

        logic [WIDTH-1:0] out_4090;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4090 (
            .a(out_4080),
            .b(out_4089),
            .outp(out_4090)
        );        
        

        logic [WIDTH-1:0] out_4091;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4091 (
            .a(out_4047),
            .b(out_4090),
            .outp(out_4091)
        );        
        

        logic [WIDTH-1:0] out_4092;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4092 (
            .in(out_4069),
            .outp(out_4092)
        );
        

        logic [WIDTH-1:0] out_4093;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.239)
        ) inst_4093 (
            .outp(out_4093)
        );
        

        logic [WIDTH-1:0] out_4094;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4094 (
            .a(out_3),
            .b(out_4093),
            .outp(out_4094)
        );        
        

        logic [WIDTH-1:0] out_4095;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4095 (
            .in(out_4094),
            .outp(out_4095)
        );
        

        logic [WIDTH-1:0] out_4096;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4096 (
            .a(out_4092),
            .b(out_4095),
            .outp(out_4096)
        );        
        

        logic [WIDTH-1:0] out_4097;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4097 (
            .in(out_4096),
            .outp(out_4097)
        );
        

        logic [WIDTH-1:0] out_4098;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4098 (
            .a(out_4097),
            .b(out_460),
            .outp(out_4098)
        );        
        

        logic [WIDTH-1:0] out_4099;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4099 (
            .a(out_4091),
            .b(out_4098),
            .outp(out_4099)
        );        
        

        logic [WIDTH-1:0] out_4100;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.781)
        ) inst_4100 (
            .outp(out_4100)
        );
        

        logic [WIDTH-1:0] out_4101;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4101 (
            .a(out_3),
            .b(out_4100),
            .outp(out_4101)
        );        
        

        logic [WIDTH-1:0] out_4102;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4102 (
            .a(out_2888),
            .b(out_4101),
            .outp(out_4102)
        );        
        

        logic [WIDTH-1:0] out_4103;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.681)
        ) inst_4103 (
            .outp(out_4103)
        );
        

        logic [WIDTH-1:0] out_4104;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4104 (
            .a(out_4103),
            .b(out_3),
            .outp(out_4104)
        );        
        

        logic [WIDTH-1:0] out_4105;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4105 (
            .a(out_4102),
            .b(out_4104),
            .outp(out_4105)
        );        
        

        logic [WIDTH-1:0] out_4106;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4106 (
            .a(out_4105),
            .b(out_2892),
            .outp(out_4106)
        );        
        

        logic [WIDTH-1:0] out_4107;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4107 (
            .a(out_4099),
            .b(out_4106),
            .outp(out_4107)
        );        
        

        logic [WIDTH-1:0] out_4108;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.23715)
        ) inst_4108 (
            .outp(out_4108)
        );
        

        logic [WIDTH-1:0] out_4109;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4109 (
            .a(out_194),
            .b(out_4108),
            .outp(out_4109)
        );        
        

        logic [WIDTH-1:0] out_4110;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4110 (
            .a(out_2888),
            .b(out_4109),
            .outp(out_4110)
        );        
        

        logic [WIDTH-1:0] out_4111;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.68715)
        ) inst_4111 (
            .outp(out_4111)
        );
        

        logic [WIDTH-1:0] out_4112;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4112 (
            .a(out_4111),
            .b(out_194),
            .outp(out_4112)
        );        
        

        logic [WIDTH-1:0] out_4113;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4113 (
            .a(out_4110),
            .b(out_4112),
            .outp(out_4113)
        );        
        

        logic [WIDTH-1:0] out_4114;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(9.04643)
        ) inst_4114 (
            .outp(out_4114)
        );
        

        logic [WIDTH-1:0] out_4115;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4115 (
            .a(out_204),
            .b(out_4114),
            .outp(out_4115)
        );        
        

        logic [WIDTH-1:0] out_4116;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4116 (
            .in(out_4115),
            .outp(out_4116)
        );
        

        logic [WIDTH-1:0] out_4117;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4117 (
            .a(out_2904),
            .b(out_4116),
            .outp(out_4117)
        );        
        

        logic [WIDTH-1:0] out_4118;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4118 (
            .in(out_4117),
            .outp(out_4118)
        );
        

        logic [WIDTH-1:0] out_4119;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4119 (
            .a(out_200),
            .b(out_4118),
            .outp(out_4119)
        );        
        

        logic [WIDTH-1:0] out_4120;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4120 (
            .a(out_4113),
            .b(out_4119),
            .outp(out_4120)
        );        
        

        logic [WIDTH-1:0] out_4121;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4121 (
            .in(out_4109),
            .outp(out_4121)
        );
        

        logic [WIDTH-1:0] out_4122;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4122 (
            .a(out_2904),
            .b(out_4121),
            .outp(out_4122)
        );        
        

        logic [WIDTH-1:0] out_4123;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4123 (
            .in(out_4122),
            .outp(out_4123)
        );
        

        logic [WIDTH-1:0] out_4124;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4124 (
            .a(out_4123),
            .b(out_214),
            .outp(out_4124)
        );        
        

        logic [WIDTH-1:0] out_4125;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4125 (
            .a(out_4120),
            .b(out_4124),
            .outp(out_4125)
        );        
        

        logic [WIDTH-1:0] out_4126;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4126 (
            .a(out_4125),
            .b(out_2892),
            .outp(out_4126)
        );        
        

        logic [WIDTH-1:0] out_4127;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4127 (
            .a(out_4107),
            .b(out_4126),
            .outp(out_4127)
        );        
        

        logic [WIDTH-1:0] out_4128;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.306)
        ) inst_4128 (
            .outp(out_4128)
        );
        

        logic [WIDTH-1:0] out_4129;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4129 (
            .a(out_3),
            .b(out_4128),
            .outp(out_4129)
        );        
        

        logic [WIDTH-1:0] out_4130;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4130 (
            .in(out_4129),
            .outp(out_4130)
        );
        

        logic [WIDTH-1:0] out_4131;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4131 (
            .a(out_2962),
            .b(out_4130),
            .outp(out_4131)
        );        
        

        logic [WIDTH-1:0] out_4132;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4132 (
            .in(out_4131),
            .outp(out_4132)
        );
        

        logic [WIDTH-1:0] out_4133;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4133 (
            .a(out_9),
            .b(out_4132),
            .outp(out_4133)
        );        
        

        logic [WIDTH-1:0] out_4134;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4134 (
            .a(out_4132),
            .b(out_21),
            .outp(out_4134)
        );        
        

        logic [WIDTH-1:0] out_4135;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4135 (
            .a(out_4133),
            .b(out_4134),
            .outp(out_4135)
        );        
        

        logic [WIDTH-1:0] out_4136;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4136 (
            .a(out_4127),
            .b(out_4135),
            .outp(out_4136)
        );        
        

        logic [WIDTH-1:0] out_4137;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.98571)
        ) inst_4137 (
            .outp(out_4137)
        );
        

        logic [WIDTH-1:0] out_4138;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4138 (
            .a(out_4137),
            .b(out_194),
            .outp(out_4138)
        );        
        

        logic [WIDTH-1:0] out_4139;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4139 (
            .a(out_1676),
            .b(out_4138),
            .outp(out_4139)
        );        
        

        logic [WIDTH-1:0] out_4140;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.53571)
        ) inst_4140 (
            .outp(out_4140)
        );
        

        logic [WIDTH-1:0] out_4141;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4141 (
            .a(out_4140),
            .b(out_194),
            .outp(out_4141)
        );        
        

        logic [WIDTH-1:0] out_4142;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4142 (
            .in(out_4141),
            .outp(out_4142)
        );
        

        logic [WIDTH-1:0] out_4143;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4143 (
            .a(out_4139),
            .b(out_4142),
            .outp(out_4143)
        );        
        

        logic [WIDTH-1:0] out_4144;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(9.98214)
        ) inst_4144 (
            .outp(out_4144)
        );
        

        logic [WIDTH-1:0] out_4145;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4145 (
            .a(out_4144),
            .b(out_204),
            .outp(out_4145)
        );        
        

        logic [WIDTH-1:0] out_4146;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4146 (
            .in(out_4145),
            .outp(out_4146)
        );
        

        logic [WIDTH-1:0] out_4147;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4147 (
            .a(out_2020),
            .b(out_4146),
            .outp(out_4147)
        );        
        

        logic [WIDTH-1:0] out_4148;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4148 (
            .in(out_4147),
            .outp(out_4148)
        );
        

        logic [WIDTH-1:0] out_4149;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4149 (
            .a(out_200),
            .b(out_4148),
            .outp(out_4149)
        );        
        

        logic [WIDTH-1:0] out_4150;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4150 (
            .a(out_4143),
            .b(out_4149),
            .outp(out_4150)
        );        
        

        logic [WIDTH-1:0] out_4151;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4151 (
            .in(out_4138),
            .outp(out_4151)
        );
        

        logic [WIDTH-1:0] out_4152;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4152 (
            .a(out_2020),
            .b(out_4151),
            .outp(out_4152)
        );        
        

        logic [WIDTH-1:0] out_4153;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4153 (
            .in(out_4152),
            .outp(out_4153)
        );
        

        logic [WIDTH-1:0] out_4154;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4154 (
            .a(out_4153),
            .b(out_214),
            .outp(out_4154)
        );        
        

        logic [WIDTH-1:0] out_4155;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4155 (
            .a(out_4150),
            .b(out_4154),
            .outp(out_4155)
        );        
        

        logic [WIDTH-1:0] out_4156;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4156 (
            .a(out_4136),
            .b(out_4155),
            .outp(out_4156)
        );        
        

        logic [WIDTH-1:0] out_4157;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.5)
        ) inst_4157 (
            .outp(out_4157)
        );
        

        logic [WIDTH-1:0] out_4158;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4158 (
            .a(out_4157),
            .b(out_3),
            .outp(out_4158)
        );        
        

        logic [WIDTH-1:0] out_4159;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4159 (
            .a(out_1870),
            .b(out_4158),
            .outp(out_4159)
        );        
        

        logic [WIDTH-1:0] out_4160;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.6)
        ) inst_4160 (
            .outp(out_4160)
        );
        

        logic [WIDTH-1:0] out_4161;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4161 (
            .a(out_4160),
            .b(out_3),
            .outp(out_4161)
        );        
        

        logic [WIDTH-1:0] out_4162;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4162 (
            .in(out_4161),
            .outp(out_4162)
        );
        

        logic [WIDTH-1:0] out_4163;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4163 (
            .a(out_4159),
            .b(out_4162),
            .outp(out_4163)
        );        
        

        logic [WIDTH-1:0] out_4164;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4164 (
            .a(out_4156),
            .b(out_4163),
            .outp(out_4164)
        );        
        

        logic [WIDTH-1:0] out_4165;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4165 (
            .a(out_1675),
            .b(out_1850),
            .outp(out_4165)
        );        
        

        logic [WIDTH-1:0] out_4166;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4166 (
            .a(out_4165),
            .b(out_1970),
            .outp(out_4166)
        );        
        

        logic [WIDTH-1:0] out_4167;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4167 (
            .in(out_4158),
            .outp(out_4167)
        );
        

        logic [WIDTH-1:0] out_4168;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4168 (
            .a(out_4166),
            .b(out_4167),
            .outp(out_4168)
        );        
        

        logic [WIDTH-1:0] out_4169;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4169 (
            .a(out_4164),
            .b(out_4168),
            .outp(out_4169)
        );        
        

        logic [WIDTH-1:0] out_4170;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4170 (
            .a(out_1660),
            .b(out_1850),
            .outp(out_4170)
        );        
        

        logic [WIDTH-1:0] out_4171;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4171 (
            .a(out_4170),
            .b(out_2081),
            .outp(out_4171)
        );        
        

        logic [WIDTH-1:0] out_4172;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4172 (
            .a(out_4171),
            .b(out_4167),
            .outp(out_4172)
        );        
        

        logic [WIDTH-1:0] out_4173;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4173 (
            .a(out_4169),
            .b(out_4172),
            .outp(out_4173)
        );        
        

        logic [WIDTH-1:0] out_4174;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.6)
        ) inst_4174 (
            .outp(out_4174)
        );
        

        logic [WIDTH-1:0] out_4175;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4175 (
            .a(out_4174),
            .b(out_3),
            .outp(out_4175)
        );        
        

        logic [WIDTH-1:0] out_4176;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4176 (
            .a(out_1870),
            .b(out_4175),
            .outp(out_4176)
        );        
        

        logic [WIDTH-1:0] out_4177;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4177 (
            .in(out_1850),
            .outp(out_4177)
        );
        

        logic [WIDTH-1:0] out_4178;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4178 (
            .a(out_4176),
            .b(out_4177),
            .outp(out_4178)
        );        
        

        logic [WIDTH-1:0] out_4179;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4179 (
            .a(out_1851),
            .b(out_1873),
            .outp(out_4179)
        );        
        

        logic [WIDTH-1:0] out_4180;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4180 (
            .in(out_4179),
            .outp(out_4180)
        );
        

        logic [WIDTH-1:0] out_4181;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4181 (
            .a(out_9),
            .b(out_4180),
            .outp(out_4181)
        );        
        

        logic [WIDTH-1:0] out_4182;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4182 (
            .a(out_4178),
            .b(out_4181),
            .outp(out_4182)
        );        
        

        logic [WIDTH-1:0] out_4183;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4183 (
            .a(out_4180),
            .b(out_21),
            .outp(out_4183)
        );        
        

        logic [WIDTH-1:0] out_4184;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4184 (
            .a(out_4182),
            .b(out_4183),
            .outp(out_4184)
        );        
        

        logic [WIDTH-1:0] out_4185;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4185 (
            .a(out_4173),
            .b(out_4184),
            .outp(out_4185)
        );        
        

        logic [WIDTH-1:0] out_4186;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4186 (
            .a(out_2985),
            .b(out_2892),
            .outp(out_4186)
        );        
        

        logic [WIDTH-1:0] out_4187;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.28901)
        ) inst_4187 (
            .outp(out_4187)
        );
        

        logic [WIDTH-1:0] out_4188;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4188 (
            .a(out_3),
            .b(out_4187),
            .outp(out_4188)
        );        
        

        logic [WIDTH-1:0] out_4189;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4189 (
            .a(out_4186),
            .b(out_4188),
            .outp(out_4189)
        );        
        

        logic [WIDTH-1:0] out_4190;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.18901)
        ) inst_4190 (
            .outp(out_4190)
        );
        

        logic [WIDTH-1:0] out_4191;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4191 (
            .a(out_4190),
            .b(out_3),
            .outp(out_4191)
        );        
        

        logic [WIDTH-1:0] out_4192;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4192 (
            .a(out_4189),
            .b(out_4191),
            .outp(out_4192)
        );        
        

        logic [WIDTH-1:0] out_4193;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4193 (
            .a(out_4185),
            .b(out_4192),
            .outp(out_4193)
        );        
        

        logic [WIDTH-1:0] out_4194;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.03901)
        ) inst_4194 (
            .outp(out_4194)
        );
        

        logic [WIDTH-1:0] out_4195;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4195 (
            .a(out_3),
            .b(out_4194),
            .outp(out_4195)
        );        
        

        logic [WIDTH-1:0] out_4196;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4196 (
            .a(out_4186),
            .b(out_4195),
            .outp(out_4196)
        );        
        

        logic [WIDTH-1:0] out_4197;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.93901)
        ) inst_4197 (
            .outp(out_4197)
        );
        

        logic [WIDTH-1:0] out_4198;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4198 (
            .a(out_4197),
            .b(out_3),
            .outp(out_4198)
        );        
        

        logic [WIDTH-1:0] out_4199;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4199 (
            .a(out_4196),
            .b(out_4198),
            .outp(out_4199)
        );        
        

        logic [WIDTH-1:0] out_4200;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4200 (
            .a(out_4193),
            .b(out_4199),
            .outp(out_4200)
        );        
        

        logic [WIDTH-1:0] out_4201;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.76837e-07)
        ) inst_4201 (
            .outp(out_4201)
        );
        

        logic [WIDTH-1:0] out_4202;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4202 (
            .a(out_14),
            .b(out_4201),
            .outp(out_4202)
        );        
        

        logic [WIDTH-1:0] out_4203;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4203 (
            .a(out_4202),
            .b(out_3078),
            .outp(out_4203)
        );        
        

        logic [WIDTH-1:0] out_4204;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.81401)
        ) inst_4204 (
            .outp(out_4204)
        );
        

        logic [WIDTH-1:0] out_4205;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4205 (
            .a(out_3),
            .b(out_4204),
            .outp(out_4205)
        );        
        

        logic [WIDTH-1:0] out_4206;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4206 (
            .a(out_4203),
            .b(out_4205),
            .outp(out_4206)
        );        
        

        logic [WIDTH-1:0] out_4207;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.71401)
        ) inst_4207 (
            .outp(out_4207)
        );
        

        logic [WIDTH-1:0] out_4208;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4208 (
            .a(out_4207),
            .b(out_3),
            .outp(out_4208)
        );        
        

        logic [WIDTH-1:0] out_4209;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4209 (
            .a(out_4206),
            .b(out_4208),
            .outp(out_4209)
        );        
        

        logic [WIDTH-1:0] out_4210;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4210 (
            .a(out_4200),
            .b(out_4209),
            .outp(out_4210)
        );        
        

        logic [WIDTH-1:0] out_4211;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.1)
        ) inst_4211 (
            .outp(out_4211)
        );
        

        logic [WIDTH-1:0] out_4212;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4212 (
            .a(out_4211),
            .b(out_14),
            .outp(out_4212)
        );        
        

        logic [WIDTH-1:0] out_4213;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4213 (
            .a(out_2985),
            .b(out_4212),
            .outp(out_4213)
        );        
        

        logic [WIDTH-1:0] out_4214;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.61401)
        ) inst_4214 (
            .outp(out_4214)
        );
        

        logic [WIDTH-1:0] out_4215;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4215 (
            .a(out_3),
            .b(out_4214),
            .outp(out_4215)
        );        
        

        logic [WIDTH-1:0] out_4216;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4216 (
            .a(out_4213),
            .b(out_4215),
            .outp(out_4216)
        );        
        

        logic [WIDTH-1:0] out_4217;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.11401)
        ) inst_4217 (
            .outp(out_4217)
        );
        

        logic [WIDTH-1:0] out_4218;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4218 (
            .a(out_4217),
            .b(out_3),
            .outp(out_4218)
        );        
        

        logic [WIDTH-1:0] out_4219;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4219 (
            .a(out_4216),
            .b(out_4218),
            .outp(out_4219)
        );        
        

        logic [WIDTH-1:0] out_4220;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4220 (
            .a(out_4210),
            .b(out_4219),
            .outp(out_4220)
        );        
        

        logic [WIDTH-1:0] out_4221;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4221 (
            .a(out_2892),
            .b(out_4215),
            .outp(out_4221)
        );        
        

        logic [WIDTH-1:0] out_4222;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4222 (
            .a(out_4221),
            .b(out_4218),
            .outp(out_4222)
        );        
        

        logic [WIDTH-1:0] out_4223;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.7)
        ) inst_4223 (
            .outp(out_4223)
        );
        

        logic [WIDTH-1:0] out_4224;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4224 (
            .a(out_4223),
            .b(out_14),
            .outp(out_4224)
        );        
        

        logic [WIDTH-1:0] out_4225;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4225 (
            .a(out_4222),
            .b(out_4224),
            .outp(out_4225)
        );        
        

        logic [WIDTH-1:0] out_4226;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4226 (
            .a(out_4220),
            .b(out_4225),
            .outp(out_4226)
        );        
        

        logic [WIDTH-1:0] out_4227;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.41401)
        ) inst_4227 (
            .outp(out_4227)
        );
        

        logic [WIDTH-1:0] out_4228;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4228 (
            .a(out_3),
            .b(out_4227),
            .outp(out_4228)
        );        
        

        logic [WIDTH-1:0] out_4229;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4229 (
            .a(out_4186),
            .b(out_4228),
            .outp(out_4229)
        );        
        

        logic [WIDTH-1:0] out_4230;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.314)
        ) inst_4230 (
            .outp(out_4230)
        );
        

        logic [WIDTH-1:0] out_4231;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4231 (
            .a(out_4230),
            .b(out_3),
            .outp(out_4231)
        );        
        

        logic [WIDTH-1:0] out_4232;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4232 (
            .a(out_4229),
            .b(out_4231),
            .outp(out_4232)
        );        
        

        logic [WIDTH-1:0] out_4233;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4233 (
            .a(out_4226),
            .b(out_4232),
            .outp(out_4233)
        );        
        

        logic [WIDTH-1:0] out_4234;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4234 (
            .a(out_2888),
            .b(out_2892),
            .outp(out_4234)
        );        
        

        logic [WIDTH-1:0] out_4235;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.1185)
        ) inst_4235 (
            .outp(out_4235)
        );
        

        logic [WIDTH-1:0] out_4236;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4236 (
            .a(out_3),
            .b(out_4235),
            .outp(out_4236)
        );        
        

        logic [WIDTH-1:0] out_4237;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4237 (
            .a(out_4234),
            .b(out_4236),
            .outp(out_4237)
        );        
        

        logic [WIDTH-1:0] out_4238;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0185)
        ) inst_4238 (
            .outp(out_4238)
        );
        

        logic [WIDTH-1:0] out_4239;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4239 (
            .a(out_4238),
            .b(out_3),
            .outp(out_4239)
        );        
        

        logic [WIDTH-1:0] out_4240;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4240 (
            .a(out_4237),
            .b(out_4239),
            .outp(out_4240)
        );        
        

        logic [WIDTH-1:0] out_4241;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4241 (
            .a(out_4233),
            .b(out_4240),
            .outp(out_4241)
        );        
        

        logic [WIDTH-1:0] out_4242;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0685)
        ) inst_4242 (
            .outp(out_4242)
        );
        

        logic [WIDTH-1:0] out_4243;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4243 (
            .a(out_3),
            .b(out_4242),
            .outp(out_4243)
        );        
        

        logic [WIDTH-1:0] out_4244;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4244 (
            .in(out_4243),
            .outp(out_4244)
        );
        

        logic [WIDTH-1:0] out_4245;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4245 (
            .a(out_2931),
            .b(out_4244),
            .outp(out_4245)
        );        
        

        logic [WIDTH-1:0] out_4246;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4246 (
            .in(out_4245),
            .outp(out_4246)
        );
        

        logic [WIDTH-1:0] out_4247;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4247 (
            .a(out_4246),
            .b(out_460),
            .outp(out_4247)
        );        
        

        logic [WIDTH-1:0] out_4248;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4248 (
            .a(out_4241),
            .b(out_4247),
            .outp(out_4248)
        );        
        

        logic [WIDTH-1:0] out_4249;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4249 (
            .a(out_2892),
            .b(out_2944),
            .outp(out_4249)
        );        
        

        logic [WIDTH-1:0] out_4250;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.1935)
        ) inst_4250 (
            .outp(out_4250)
        );
        

        logic [WIDTH-1:0] out_4251;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4251 (
            .a(out_3),
            .b(out_4250),
            .outp(out_4251)
        );        
        

        logic [WIDTH-1:0] out_4252;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4252 (
            .a(out_4249),
            .b(out_4251),
            .outp(out_4252)
        );        
        

        logic [WIDTH-1:0] out_4253;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.0935)
        ) inst_4253 (
            .outp(out_4253)
        );
        

        logic [WIDTH-1:0] out_4254;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4254 (
            .a(out_4253),
            .b(out_3),
            .outp(out_4254)
        );        
        

        logic [WIDTH-1:0] out_4255;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4255 (
            .a(out_4252),
            .b(out_4254),
            .outp(out_4255)
        );        
        

        logic [WIDTH-1:0] out_4256;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4256 (
            .a(out_4248),
            .b(out_4255),
            .outp(out_4256)
        );        
        

        logic [WIDTH-1:0] out_4257;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.943501)
        ) inst_4257 (
            .outp(out_4257)
        );
        

        logic [WIDTH-1:0] out_4258;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4258 (
            .a(out_3),
            .b(out_4257),
            .outp(out_4258)
        );        
        

        logic [WIDTH-1:0] out_4259;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4259 (
            .a(out_4249),
            .b(out_4258),
            .outp(out_4259)
        );        
        

        logic [WIDTH-1:0] out_4260;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.8435)
        ) inst_4260 (
            .outp(out_4260)
        );
        

        logic [WIDTH-1:0] out_4261;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4261 (
            .a(out_4260),
            .b(out_3),
            .outp(out_4261)
        );        
        

        logic [WIDTH-1:0] out_4262;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4262 (
            .a(out_4259),
            .b(out_4261),
            .outp(out_4262)
        );        
        

        logic [WIDTH-1:0] out_4263;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4263 (
            .a(out_4256),
            .b(out_4262),
            .outp(out_4263)
        );        
        

        logic [WIDTH-1:0] out_4264;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.275)
        ) inst_4264 (
            .outp(out_4264)
        );
        

        logic [WIDTH-1:0] out_4265;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4265 (
            .a(out_4264),
            .b(out_14),
            .outp(out_4265)
        );        
        

        logic [WIDTH-1:0] out_4266;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4266 (
            .a(out_2892),
            .b(out_4265),
            .outp(out_4266)
        );        
        

        logic [WIDTH-1:0] out_4267;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.693501)
        ) inst_4267 (
            .outp(out_4267)
        );
        

        logic [WIDTH-1:0] out_4268;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4268 (
            .a(out_3),
            .b(out_4267),
            .outp(out_4268)
        );        
        

        logic [WIDTH-1:0] out_4269;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4269 (
            .a(out_4266),
            .b(out_4268),
            .outp(out_4269)
        );        
        

        logic [WIDTH-1:0] out_4270;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5935)
        ) inst_4270 (
            .outp(out_4270)
        );
        

        logic [WIDTH-1:0] out_4271;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4271 (
            .a(out_4270),
            .b(out_3),
            .outp(out_4271)
        );        
        

        logic [WIDTH-1:0] out_4272;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4272 (
            .a(out_4269),
            .b(out_4271),
            .outp(out_4272)
        );        
        

        logic [WIDTH-1:0] out_4273;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4273 (
            .a(out_4263),
            .b(out_4272),
            .outp(out_4273)
        );        
        

        logic [WIDTH-1:0] out_4274;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4274 (
            .a(out_4271),
            .b(out_3081),
            .outp(out_4274)
        );        
        

        logic [WIDTH-1:0] out_4275;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.45)
        ) inst_4275 (
            .outp(out_4275)
        );
        

        logic [WIDTH-1:0] out_4276;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4276 (
            .a(out_4275),
            .b(out_14),
            .outp(out_4276)
        );        
        

        logic [WIDTH-1:0] out_4277;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4277 (
            .in(out_4276),
            .outp(out_4277)
        );
        

        logic [WIDTH-1:0] out_4278;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4278 (
            .a(out_4274),
            .b(out_4277),
            .outp(out_4278)
        );        
        

        logic [WIDTH-1:0] out_4279;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2435)
        ) inst_4279 (
            .outp(out_4279)
        );
        

        logic [WIDTH-1:0] out_4280;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4280 (
            .a(out_3),
            .b(out_4279),
            .outp(out_4280)
        );        
        

        logic [WIDTH-1:0] out_4281;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4281 (
            .a(out_4278),
            .b(out_4280),
            .outp(out_4281)
        );        
        

        logic [WIDTH-1:0] out_4282;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4282 (
            .in(out_2944),
            .outp(out_4282)
        );
        

        logic [WIDTH-1:0] out_4283;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.0185)
        ) inst_4283 (
            .outp(out_4283)
        );
        

        logic [WIDTH-1:0] out_4284;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4284 (
            .a(out_3),
            .b(out_4283),
            .outp(out_4284)
        );        
        

        logic [WIDTH-1:0] out_4285;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4285 (
            .in(out_4284),
            .outp(out_4285)
        );
        

        logic [WIDTH-1:0] out_4286;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4286 (
            .a(out_4282),
            .b(out_4285),
            .outp(out_4286)
        );        
        

        logic [WIDTH-1:0] out_4287;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4287 (
            .in(out_4286),
            .outp(out_4287)
        );
        

        logic [WIDTH-1:0] out_4288;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4288 (
            .a(out_460),
            .b(out_4287),
            .outp(out_4288)
        );        
        

        logic [WIDTH-1:0] out_4289;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4289 (
            .a(out_4287),
            .b(out_9),
            .outp(out_4289)
        );        
        

        logic [WIDTH-1:0] out_4290;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4290 (
            .a(out_4288),
            .b(out_4289),
            .outp(out_4290)
        );        
        

        logic [WIDTH-1:0] out_4291;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.7685)
        ) inst_4291 (
            .outp(out_4291)
        );
        

        logic [WIDTH-1:0] out_4292;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4292 (
            .a(out_3),
            .b(out_4291),
            .outp(out_4292)
        );        
        

        logic [WIDTH-1:0] out_4293;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4293 (
            .in(out_4292),
            .outp(out_4293)
        );
        

        logic [WIDTH-1:0] out_4294;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4294 (
            .a(out_4282),
            .b(out_4293),
            .outp(out_4294)
        );        
        

        logic [WIDTH-1:0] out_4295;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4295 (
            .in(out_4294),
            .outp(out_4295)
        );
        

        logic [WIDTH-1:0] out_4296;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4296 (
            .a(out_460),
            .b(out_4295),
            .outp(out_4296)
        );        
        

        logic [WIDTH-1:0] out_4297;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4297 (
            .a(out_4295),
            .b(out_9),
            .outp(out_4297)
        );        
        

        logic [WIDTH-1:0] out_4298;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4298 (
            .a(out_4296),
            .b(out_4297),
            .outp(out_4298)
        );        
        

        logic [WIDTH-1:0] out_4299;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4299 (
            .a(out_4290),
            .b(out_4298),
            .outp(out_4299)
        );        
        

        logic [WIDTH-1:0] out_4300;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4300 (
            .a(out_4281),
            .b(out_4299),
            .outp(out_4300)
        );        
        

        logic [WIDTH-1:0] out_4301;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4301 (
            .a(out_4273),
            .b(out_4300),
            .outp(out_4301)
        );        
        

        logic [WIDTH-1:0] out_4302;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.2355)
        ) inst_4302 (
            .outp(out_4302)
        );
        

        logic [WIDTH-1:0] out_4303;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4303 (
            .a(out_3),
            .b(out_4302),
            .outp(out_4303)
        );        
        

        logic [WIDTH-1:0] out_4304;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4304 (
            .a(out_4234),
            .b(out_4303),
            .outp(out_4304)
        );        
        

        logic [WIDTH-1:0] out_4305;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.1355)
        ) inst_4305 (
            .outp(out_4305)
        );
        

        logic [WIDTH-1:0] out_4306;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4306 (
            .a(out_4305),
            .b(out_3),
            .outp(out_4306)
        );        
        

        logic [WIDTH-1:0] out_4307;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4307 (
            .a(out_4304),
            .b(out_4306),
            .outp(out_4307)
        );        
        

        logic [WIDTH-1:0] out_4308;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4308 (
            .a(out_4301),
            .b(out_4307),
            .outp(out_4308)
        );        
        

        logic [WIDTH-1:0] out_4309;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0499997)
        ) inst_4309 (
            .outp(out_4309)
        );
        

        logic [WIDTH-1:0] out_4310;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4310 (
            .a(out_4309),
            .b(out_14),
            .outp(out_4310)
        );        
        

        logic [WIDTH-1:0] out_4311;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.781)
        ) inst_4311 (
            .outp(out_4311)
        );
        

        logic [WIDTH-1:0] out_4312;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4312 (
            .a(out_3),
            .b(out_4311),
            .outp(out_4312)
        );        
        

        logic [WIDTH-1:0] out_4313;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4313 (
            .a(out_4310),
            .b(out_4312),
            .outp(out_4313)
        );        
        

        logic [WIDTH-1:0] out_4314;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4314 (
            .a(out_4313),
            .b(out_2892),
            .outp(out_4314)
        );        
        

        logic [WIDTH-1:0] out_4315;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.681)
        ) inst_4315 (
            .outp(out_4315)
        );
        

        logic [WIDTH-1:0] out_4316;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4316 (
            .a(out_4315),
            .b(out_3),
            .outp(out_4316)
        );        
        

        logic [WIDTH-1:0] out_4317;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4317 (
            .a(out_4314),
            .b(out_4316),
            .outp(out_4317)
        );        
        

        logic [WIDTH-1:0] out_4318;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4318 (
            .a(out_4308),
            .b(out_4317),
            .outp(out_4318)
        );        
        

        logic [WIDTH-1:0] out_4319;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.35)
        ) inst_4319 (
            .outp(out_4319)
        );
        

        logic [WIDTH-1:0] out_4320;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4320 (
            .a(out_4319),
            .b(out_14),
            .outp(out_4320)
        );        
        

        logic [WIDTH-1:0] out_4321;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4321 (
            .in(out_4320),
            .outp(out_4321)
        );
        

        logic [WIDTH-1:0] out_4322;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4322 (
            .a(out_2888),
            .b(out_4321),
            .outp(out_4322)
        );        
        

        logic [WIDTH-1:0] out_4323;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.931)
        ) inst_4323 (
            .outp(out_4323)
        );
        

        logic [WIDTH-1:0] out_4324;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4324 (
            .a(out_3),
            .b(out_4323),
            .outp(out_4324)
        );        
        

        logic [WIDTH-1:0] out_4325;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4325 (
            .a(out_4322),
            .b(out_4324),
            .outp(out_4325)
        );        
        

        logic [WIDTH-1:0] out_4326;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.531)
        ) inst_4326 (
            .outp(out_4326)
        );
        

        logic [WIDTH-1:0] out_4327;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4327 (
            .a(out_4326),
            .b(out_3),
            .outp(out_4327)
        );        
        

        logic [WIDTH-1:0] out_4328;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4328 (
            .a(out_4325),
            .b(out_4327),
            .outp(out_4328)
        );        
        

        logic [WIDTH-1:0] out_4329;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4329 (
            .a(out_4318),
            .b(out_4328),
            .outp(out_4329)
        );        
        

        logic [WIDTH-1:0] out_4330;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4330 (
            .a(out_2985),
            .b(out_4324),
            .outp(out_4330)
        );        
        

        logic [WIDTH-1:0] out_4331;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4331 (
            .a(out_4330),
            .b(out_4327),
            .outp(out_4331)
        );        
        

        logic [WIDTH-1:0] out_4332;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4332 (
            .in(out_4310),
            .outp(out_4332)
        );
        

        logic [WIDTH-1:0] out_4333;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4333 (
            .a(out_4331),
            .b(out_4332),
            .outp(out_4333)
        );        
        

        logic [WIDTH-1:0] out_4334;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4334 (
            .in(out_4310),
            .outp(out_4334)
        );
        

        logic [WIDTH-1:0] out_4335;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4335 (
            .in(out_4324),
            .outp(out_4335)
        );
        

        logic [WIDTH-1:0] out_4336;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4336 (
            .a(out_4334),
            .b(out_4335),
            .outp(out_4336)
        );        
        

        logic [WIDTH-1:0] out_4337;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4337 (
            .in(out_4336),
            .outp(out_4337)
        );
        

        logic [WIDTH-1:0] out_4338;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4338 (
            .a(out_336),
            .b(out_4337),
            .outp(out_4338)
        );        
        

        logic [WIDTH-1:0] out_4339;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4339 (
            .a(out_4333),
            .b(out_4338),
            .outp(out_4339)
        );        
        

        logic [WIDTH-1:0] out_4340;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4340 (
            .a(out_4337),
            .b(out_343),
            .outp(out_4340)
        );        
        

        logic [WIDTH-1:0] out_4341;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4341 (
            .a(out_4339),
            .b(out_4340),
            .outp(out_4341)
        );        
        

        logic [WIDTH-1:0] out_4342;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4342 (
            .a(out_4329),
            .b(out_4341),
            .outp(out_4342)
        );        
        

        logic [WIDTH-1:0] out_4343;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4343 (
            .a(out_3176),
            .b(out_3179),
            .outp(out_4343)
        );        
        

        logic [WIDTH-1:0] out_4344;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.65817)
        ) inst_4344 (
            .outp(out_4344)
        );
        

        logic [WIDTH-1:0] out_4345;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4345 (
            .a(out_4344),
            .b(out_260),
            .outp(out_4345)
        );        
        

        logic [WIDTH-1:0] out_4346;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4346 (
            .a(out_4343),
            .b(out_4345),
            .outp(out_4346)
        );        
        

        logic [WIDTH-1:0] out_4347;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.82067)
        ) inst_4347 (
            .outp(out_4347)
        );
        

        logic [WIDTH-1:0] out_4348;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4348 (
            .a(out_260),
            .b(out_4347),
            .outp(out_4348)
        );        
        

        logic [WIDTH-1:0] out_4349;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4349 (
            .a(out_4346),
            .b(out_4348),
            .outp(out_4349)
        );        
        

        logic [WIDTH-1:0] out_4350;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.10378)
        ) inst_4350 (
            .outp(out_4350)
        );
        

        logic [WIDTH-1:0] out_4351;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4351 (
            .a(out_4350),
            .b(out_241),
            .outp(out_4351)
        );        
        

        logic [WIDTH-1:0] out_4352;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4352 (
            .in(out_4351),
            .outp(out_4352)
        );
        

        logic [WIDTH-1:0] out_4353;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4353 (
            .a(out_3188),
            .b(out_4352),
            .outp(out_4353)
        );        
        

        logic [WIDTH-1:0] out_4354;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4354 (
            .in(out_4353),
            .outp(out_4354)
        );
        

        logic [WIDTH-1:0] out_4355;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4355 (
            .a(out_4354),
            .b(out_250),
            .outp(out_4355)
        );        
        

        logic [WIDTH-1:0] out_4356;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4356 (
            .a(out_4349),
            .b(out_4355),
            .outp(out_4356)
        );        
        

        logic [WIDTH-1:0] out_4357;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4357 (
            .in(out_4356),
            .outp(out_4357)
        );
        

        logic [WIDTH-1:0] out_4358;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4358 (
            .in(out_4345),
            .outp(out_4358)
        );
        

        logic [WIDTH-1:0] out_4359;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4359 (
            .a(out_3198),
            .b(out_4358),
            .outp(out_4359)
        );        
        

        logic [WIDTH-1:0] out_4360;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4360 (
            .in(out_4359),
            .outp(out_4360)
        );
        

        logic [WIDTH-1:0] out_4361;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4361 (
            .a(out_4360),
            .b(out_275),
            .outp(out_4361)
        );        
        

        logic [WIDTH-1:0] out_4362;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4362 (
            .a(out_4357),
            .b(out_4361),
            .outp(out_4362)
        );        
        

        logic [WIDTH-1:0] out_4363;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4363 (
            .a(out_4342),
            .b(out_4362),
            .outp(out_4363)
        );        
        

        logic [WIDTH-1:0] out_4364;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4364 (
            .a(out_3211),
            .b(out_3215),
            .outp(out_4364)
        );        
        

        logic [WIDTH-1:0] out_4365;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.65817)
        ) inst_4365 (
            .outp(out_4365)
        );
        

        logic [WIDTH-1:0] out_4366;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4366 (
            .a(out_260),
            .b(out_4365),
            .outp(out_4366)
        );        
        

        logic [WIDTH-1:0] out_4367;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4367 (
            .a(out_4364),
            .b(out_4366),
            .outp(out_4367)
        );        
        

        logic [WIDTH-1:0] out_4368;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.49567)
        ) inst_4368 (
            .outp(out_4368)
        );
        

        logic [WIDTH-1:0] out_4369;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4369 (
            .a(out_4368),
            .b(out_260),
            .outp(out_4369)
        );        
        

        logic [WIDTH-1:0] out_4370;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4370 (
            .a(out_4367),
            .b(out_4369),
            .outp(out_4370)
        );        
        

        logic [WIDTH-1:0] out_4371;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.10711)
        ) inst_4371 (
            .outp(out_4371)
        );
        

        logic [WIDTH-1:0] out_4372;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4372 (
            .a(out_241),
            .b(out_4371),
            .outp(out_4372)
        );        
        

        logic [WIDTH-1:0] out_4373;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4373 (
            .in(out_4372),
            .outp(out_4373)
        );
        

        logic [WIDTH-1:0] out_4374;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4374 (
            .a(out_3222),
            .b(out_4373),
            .outp(out_4374)
        );        
        

        logic [WIDTH-1:0] out_4375;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4375 (
            .in(out_4374),
            .outp(out_4375)
        );
        

        logic [WIDTH-1:0] out_4376;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4376 (
            .a(out_4375),
            .b(out_250),
            .outp(out_4376)
        );        
        

        logic [WIDTH-1:0] out_4377;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4377 (
            .a(out_4370),
            .b(out_4376),
            .outp(out_4377)
        );        
        

        logic [WIDTH-1:0] out_4378;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4378 (
            .in(out_4377),
            .outp(out_4378)
        );
        

        logic [WIDTH-1:0] out_4379;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4379 (
            .in(out_4366),
            .outp(out_4379)
        );
        

        logic [WIDTH-1:0] out_4380;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4380 (
            .a(out_3231),
            .b(out_4379),
            .outp(out_4380)
        );        
        

        logic [WIDTH-1:0] out_4381;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4381 (
            .in(out_4380),
            .outp(out_4381)
        );
        

        logic [WIDTH-1:0] out_4382;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4382 (
            .a(out_4381),
            .b(out_275),
            .outp(out_4382)
        );        
        

        logic [WIDTH-1:0] out_4383;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4383 (
            .a(out_4378),
            .b(out_4382),
            .outp(out_4383)
        );        
        

        logic [WIDTH-1:0] out_4384;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4384 (
            .a(out_4363),
            .b(out_4383),
            .outp(out_4384)
        );        
        

        logic [WIDTH-1:0] out_4385;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.743571)
        ) inst_4385 (
            .outp(out_4385)
        );
        

        logic [WIDTH-1:0] out_4386;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4386 (
            .a(out_194),
            .b(out_4385),
            .outp(out_4386)
        );        
        

        logic [WIDTH-1:0] out_4387;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4387 (
            .a(out_4234),
            .b(out_4386),
            .outp(out_4387)
        );        
        

        logic [WIDTH-1:0] out_4388;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.193571)
        ) inst_4388 (
            .outp(out_4388)
        );
        

        logic [WIDTH-1:0] out_4389;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4389 (
            .a(out_4388),
            .b(out_194),
            .outp(out_4389)
        );        
        

        logic [WIDTH-1:0] out_4390;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4390 (
            .a(out_4387),
            .b(out_4389),
            .outp(out_4390)
        );        
        

        logic [WIDTH-1:0] out_4391;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.929465)
        ) inst_4391 (
            .outp(out_4391)
        );
        

        logic [WIDTH-1:0] out_4392;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4392 (
            .a(out_204),
            .b(out_4391),
            .outp(out_4392)
        );        
        

        logic [WIDTH-1:0] out_4393;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4393 (
            .in(out_4392),
            .outp(out_4393)
        );
        

        logic [WIDTH-1:0] out_4394;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4394 (
            .a(out_2904),
            .b(out_4393),
            .outp(out_4394)
        );        
        

        logic [WIDTH-1:0] out_4395;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4395 (
            .in(out_4394),
            .outp(out_4395)
        );
        

        logic [WIDTH-1:0] out_4396;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4396 (
            .a(out_200),
            .b(out_4395),
            .outp(out_4396)
        );        
        

        logic [WIDTH-1:0] out_4397;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4397 (
            .a(out_4390),
            .b(out_4396),
            .outp(out_4397)
        );        
        

        logic [WIDTH-1:0] out_4398;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4398 (
            .in(out_4386),
            .outp(out_4398)
        );
        

        logic [WIDTH-1:0] out_4399;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4399 (
            .a(out_2904),
            .b(out_4398),
            .outp(out_4399)
        );        
        

        logic [WIDTH-1:0] out_4400;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4400 (
            .in(out_4399),
            .outp(out_4400)
        );
        

        logic [WIDTH-1:0] out_4401;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4401 (
            .a(out_4400),
            .b(out_214),
            .outp(out_4401)
        );        
        

        logic [WIDTH-1:0] out_4402;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4402 (
            .a(out_4397),
            .b(out_4401),
            .outp(out_4402)
        );        
        

        logic [WIDTH-1:0] out_4403;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4403 (
            .a(out_4384),
            .b(out_4402),
            .outp(out_4403)
        );        
        

        logic [WIDTH-1:0] out_4404;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(100000000.0)
        ) inst_4404 (
            .outp(out_4404)
        );
        

        logic [WIDTH-1:0] out_4405;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4405 (
            .a(out_4403),
            .b(out_4404),
            .outp(out_4405)
        );        
        

        logic [WIDTH-1:0] out_4406;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.815)
        ) inst_4406 (
            .outp(out_4406)
        );
        

        logic [WIDTH-1:0] out_4407;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4407 (
            .a(out_14),
            .b(out_4406),
            .outp(out_4407)
        );        
        

        logic [WIDTH-1:0] out_4408;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4408 (
            .a(out_1340),
            .b(out_14),
            .outp(out_4408)
        );        
        

        logic [WIDTH-1:0] out_4409;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4409 (
            .a(out_4407),
            .b(out_4408),
            .outp(out_4409)
        );        
        

        logic [WIDTH-1:0] out_4410;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.40251)
        ) inst_4410 (
            .outp(out_4410)
        );
        

        logic [WIDTH-1:0] out_4411;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4411 (
            .a(out_3),
            .b(out_4410),
            .outp(out_4411)
        );        
        

        logic [WIDTH-1:0] out_4412;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4412 (
            .a(out_4409),
            .b(out_4411),
            .outp(out_4412)
        );        
        

        logic [WIDTH-1:0] out_4413;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.90251)
        ) inst_4413 (
            .outp(out_4413)
        );
        

        logic [WIDTH-1:0] out_4414;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4414 (
            .a(out_4413),
            .b(out_3),
            .outp(out_4414)
        );        
        

        logic [WIDTH-1:0] out_4415;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4415 (
            .a(out_4412),
            .b(out_4414),
            .outp(out_4415)
        );        
        

        logic [WIDTH-1:0] out_4416;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.12751)
        ) inst_4416 (
            .outp(out_4416)
        );
        

        logic [WIDTH-1:0] out_4417;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4417 (
            .a(out_3),
            .b(out_4416),
            .outp(out_4417)
        );        
        

        logic [WIDTH-1:0] out_4418;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4418 (
            .in(out_4417),
            .outp(out_4418)
        );
        

        logic [WIDTH-1:0] out_4419;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4419 (
            .a(out_14),
            .b(out_1787),
            .outp(out_4419)
        );        
        

        logic [WIDTH-1:0] out_4420;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4420 (
            .in(out_4419),
            .outp(out_4420)
        );
        

        logic [WIDTH-1:0] out_4421;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4421 (
            .a(out_4418),
            .b(out_4420),
            .outp(out_4421)
        );        
        

        logic [WIDTH-1:0] out_4422;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4422 (
            .in(out_4421),
            .outp(out_4422)
        );
        

        logic [WIDTH-1:0] out_4423;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4423 (
            .a(out_4422),
            .b(out_21),
            .outp(out_4423)
        );        
        

        logic [WIDTH-1:0] out_4424;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.80375)
        ) inst_4424 (
            .outp(out_4424)
        );
        

        logic [WIDTH-1:0] out_4425;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4425 (
            .a(out_553),
            .b(out_4424),
            .outp(out_4425)
        );        
        

        logic [WIDTH-1:0] out_4426;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.67444)
        ) inst_4426 (
            .outp(out_4426)
        );
        

        logic [WIDTH-1:0] out_4427;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4427 (
            .a(out_559),
            .b(out_4426),
            .outp(out_4427)
        );        
        

        logic [WIDTH-1:0] out_4428;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4428 (
            .a(out_556),
            .b(out_4427),
            .outp(out_4428)
        );        
        

        logic [WIDTH-1:0] out_4429;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4429 (
            .a(out_4425),
            .b(out_4428),
            .outp(out_4429)
        );        
        

        logic [WIDTH-1:0] out_4430;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.29944)
        ) inst_4430 (
            .outp(out_4430)
        );
        

        logic [WIDTH-1:0] out_4431;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4431 (
            .a(out_4430),
            .b(out_2653),
            .outp(out_4431)
        );        
        

        logic [WIDTH-1:0] out_4432;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4432 (
            .a(out_4429),
            .b(out_4431),
            .outp(out_4432)
        );        
        

        logic [WIDTH-1:0] out_4433;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4433 (
            .a(out_2653),
            .b(out_4430),
            .outp(out_4433)
        );        
        

        logic [WIDTH-1:0] out_4434;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4434 (
            .a(out_4427),
            .b(out_556),
            .outp(out_4434)
        );        
        

        logic [WIDTH-1:0] out_4435;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4435 (
            .a(out_4433),
            .b(out_4434),
            .outp(out_4435)
        );        
        

        logic [WIDTH-1:0] out_4436;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4436 (
            .a(out_4424),
            .b(out_553),
            .outp(out_4436)
        );        
        

        logic [WIDTH-1:0] out_4437;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4437 (
            .a(out_4435),
            .b(out_4436),
            .outp(out_4437)
        );        
        

        logic [WIDTH-1:0] out_4438;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4438 (
            .a(out_4432),
            .b(out_4437),
            .outp(out_4438)
        );        
        

        logic [WIDTH-1:0] out_4439;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4439 (
            .in(out_4438),
            .outp(out_4439)
        );
        

        logic [WIDTH-1:0] out_4440;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4440 (
            .a(out_4423),
            .b(out_4439),
            .outp(out_4440)
        );        
        

        logic [WIDTH-1:0] out_4441;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4441 (
            .a(out_9),
            .b(out_4422),
            .outp(out_4441)
        );        
        

        logic [WIDTH-1:0] out_4442;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4442 (
            .a(out_4440),
            .b(out_4441),
            .outp(out_4442)
        );        
        

        logic [WIDTH-1:0] out_4443;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4443 (
            .a(out_4415),
            .b(out_4442),
            .outp(out_4443)
        );        
        

        logic [WIDTH-1:0] out_4444;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4444 (
            .a(out_4423),
            .b(out_4443),
            .outp(out_4444)
        );        
        

        logic [WIDTH-1:0] out_4445;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4445 (
            .a(out_4405),
            .b(out_4444),
            .outp(out_4445)
        );        
        

        logic [WIDTH-1:0] out_4446;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.25)
        ) inst_4446 (
            .outp(out_4446)
        );
        

        logic [WIDTH-1:0] out_4447;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4447 (
            .a(out_4446),
            .b(out_152),
            .outp(out_4447)
        );        
        

        logic [WIDTH-1:0] out_4448;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.95138)
        ) inst_4448 (
            .outp(out_4448)
        );
        

        logic [WIDTH-1:0] out_4449;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4449 (
            .a(out_131),
            .b(out_4448),
            .outp(out_4449)
        );        
        

        logic [WIDTH-1:0] out_4450;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4450 (
            .a(out_127),
            .b(out_4449),
            .outp(out_4450)
        );        
        

        logic [WIDTH-1:0] out_4451;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4451 (
            .a(out_4447),
            .b(out_4450),
            .outp(out_4451)
        );        
        

        logic [WIDTH-1:0] out_4452;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.64638)
        ) inst_4452 (
            .outp(out_4452)
        );
        

        logic [WIDTH-1:0] out_4453;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4453 (
            .a(out_4452),
            .b(out_124),
            .outp(out_4453)
        );        
        

        logic [WIDTH-1:0] out_4454;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4454 (
            .a(out_4453),
            .b(out_127),
            .outp(out_4454)
        );        
        

        logic [WIDTH-1:0] out_4455;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4455 (
            .a(out_4451),
            .b(out_4454),
            .outp(out_4455)
        );        
        

        logic [WIDTH-1:0] out_4456;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4456 (
            .a(out_4445),
            .b(out_4455),
            .outp(out_4456)
        );        
        

        logic [WIDTH-1:0] out_4457;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4457 (
            .a(out_127),
            .b(out_4453),
            .outp(out_4457)
        );        
        

        logic [WIDTH-1:0] out_4458;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4458 (
            .a(out_4449),
            .b(out_127),
            .outp(out_4458)
        );        
        

        logic [WIDTH-1:0] out_4459;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4459 (
            .a(out_4457),
            .b(out_4458),
            .outp(out_4459)
        );        
        

        logic [WIDTH-1:0] out_4460;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4460 (
            .a(out_152),
            .b(out_4446),
            .outp(out_4460)
        );        
        

        logic [WIDTH-1:0] out_4461;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4461 (
            .a(out_4459),
            .b(out_4460),
            .outp(out_4461)
        );        
        

        logic [WIDTH-1:0] out_4462;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4462 (
            .a(out_4456),
            .b(out_4461),
            .outp(out_4462)
        );        
        

        logic [WIDTH-1:0] out_4463;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.305)
        ) inst_4463 (
            .outp(out_4463)
        );
        

        logic [WIDTH-1:0] out_4464;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4464 (
            .a(out_137),
            .b(out_4463),
            .outp(out_4464)
        );        
        

        logic [WIDTH-1:0] out_4465;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4465 (
            .a(out_4457),
            .b(out_4464),
            .outp(out_4465)
        );        
        

        logic [WIDTH-1:0] out_4466;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.89638)
        ) inst_4466 (
            .outp(out_4466)
        );
        

        logic [WIDTH-1:0] out_4467;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4467 (
            .a(out_131),
            .b(out_4466),
            .outp(out_4467)
        );        
        

        logic [WIDTH-1:0] out_4468;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4468 (
            .a(out_4467),
            .b(out_127),
            .outp(out_4468)
        );        
        

        logic [WIDTH-1:0] out_4469;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4469 (
            .a(out_4465),
            .b(out_4468),
            .outp(out_4469)
        );        
        

        logic [WIDTH-1:0] out_4470;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4470 (
            .a(out_4462),
            .b(out_4469),
            .outp(out_4470)
        );        
        

        logic [WIDTH-1:0] out_4471;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4471 (
            .a(out_127),
            .b(out_4467),
            .outp(out_4471)
        );        
        

        logic [WIDTH-1:0] out_4472;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4472 (
            .a(out_4454),
            .b(out_4471),
            .outp(out_4472)
        );        
        

        logic [WIDTH-1:0] out_4473;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4473 (
            .a(out_4463),
            .b(out_137),
            .outp(out_4473)
        );        
        

        logic [WIDTH-1:0] out_4474;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4474 (
            .a(out_4472),
            .b(out_4473),
            .outp(out_4474)
        );        
        

        logic [WIDTH-1:0] out_4475;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4475 (
            .a(out_4470),
            .b(out_4474),
            .outp(out_4475)
        );        
        

        logic [WIDTH-1:0] out_4476;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.14638)
        ) inst_4476 (
            .outp(out_4476)
        );
        

        logic [WIDTH-1:0] out_4477;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4477 (
            .a(out_131),
            .b(out_127),
            .outp(out_4477)
        );        
        

        logic [WIDTH-1:0] out_4478;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4478 (
            .a(out_4476),
            .b(out_4477),
            .outp(out_4478)
        );        
        

        logic [WIDTH-1:0] out_4479;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4479 (
            .a(out_4447),
            .b(out_4478),
            .outp(out_4479)
        );        
        

        logic [WIDTH-1:0] out_4480;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4480 (
            .a(out_124),
            .b(out_127),
            .outp(out_4480)
        );        
        

        logic [WIDTH-1:0] out_4481;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.45138)
        ) inst_4481 (
            .outp(out_4481)
        );
        

        logic [WIDTH-1:0] out_4482;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4482 (
            .a(out_4480),
            .b(out_4481),
            .outp(out_4482)
        );        
        

        logic [WIDTH-1:0] out_4483;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4483 (
            .a(out_4479),
            .b(out_4482),
            .outp(out_4483)
        );        
        

        logic [WIDTH-1:0] out_4484;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4484 (
            .a(out_4475),
            .b(out_4483),
            .outp(out_4484)
        );        
        

        logic [WIDTH-1:0] out_4485;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4485 (
            .a(out_4481),
            .b(out_4480),
            .outp(out_4485)
        );        
        

        logic [WIDTH-1:0] out_4486;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4486 (
            .a(out_4460),
            .b(out_4485),
            .outp(out_4486)
        );        
        

        logic [WIDTH-1:0] out_4487;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4487 (
            .a(out_4477),
            .b(out_4476),
            .outp(out_4487)
        );        
        

        logic [WIDTH-1:0] out_4488;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4488 (
            .a(out_4486),
            .b(out_4487),
            .outp(out_4488)
        );        
        

        logic [WIDTH-1:0] out_4489;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4489 (
            .a(out_4484),
            .b(out_4488),
            .outp(out_4489)
        );        
        

        logic [WIDTH-1:0] out_4490;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4490 (
            .a(out_4464),
            .b(out_4485),
            .outp(out_4490)
        );        
        

        logic [WIDTH-1:0] out_4491;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.20138)
        ) inst_4491 (
            .outp(out_4491)
        );
        

        logic [WIDTH-1:0] out_4492;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4492 (
            .a(out_4477),
            .b(out_4491),
            .outp(out_4492)
        );        
        

        logic [WIDTH-1:0] out_4493;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4493 (
            .a(out_4490),
            .b(out_4492),
            .outp(out_4493)
        );        
        

        logic [WIDTH-1:0] out_4494;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4494 (
            .a(out_4489),
            .b(out_4493),
            .outp(out_4494)
        );        
        

        logic [WIDTH-1:0] out_4495;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4495 (
            .a(out_4473),
            .b(out_4482),
            .outp(out_4495)
        );        
        

        logic [WIDTH-1:0] out_4496;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4496 (
            .a(out_4491),
            .b(out_4477),
            .outp(out_4496)
        );        
        

        logic [WIDTH-1:0] out_4497;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4497 (
            .a(out_4495),
            .b(out_4496),
            .outp(out_4497)
        );        
        

        logic [WIDTH-1:0] out_4498;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4498 (
            .a(out_4494),
            .b(out_4497),
            .outp(out_4498)
        );        
        

        logic [WIDTH-1:0] out_4499;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8125)
        ) inst_4499 (
            .outp(out_4499)
        );
        

        logic [WIDTH-1:0] out_4500;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4500 (
            .a(out_131),
            .b(out_4499),
            .outp(out_4500)
        );        
        

        logic [WIDTH-1:0] out_4501;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4501 (
            .a(out_4500),
            .b(out_127),
            .outp(out_4501)
        );        
        

        logic [WIDTH-1:0] out_4502;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4502 (
            .in(out_4501),
            .outp(out_4502)
        );
        

        logic [WIDTH-1:0] out_4503;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6175)
        ) inst_4503 (
            .outp(out_4503)
        );
        

        logic [WIDTH-1:0] out_4504;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4504 (
            .a(out_4503),
            .b(out_124),
            .outp(out_4504)
        );        
        

        logic [WIDTH-1:0] out_4505;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4505 (
            .a(out_4504),
            .b(out_127),
            .outp(out_4505)
        );        
        

        logic [WIDTH-1:0] out_4506;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4506 (
            .a(out_4502),
            .b(out_4505),
            .outp(out_4506)
        );        
        

        logic [WIDTH-1:0] out_4507;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.14)
        ) inst_4507 (
            .outp(out_4507)
        );
        

        logic [WIDTH-1:0] out_4508;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4508 (
            .a(out_4507),
            .b(out_152),
            .outp(out_4508)
        );        
        

        logic [WIDTH-1:0] out_4509;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4509 (
            .a(out_4506),
            .b(out_4508),
            .outp(out_4509)
        );        
        

        logic [WIDTH-1:0] out_4510;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4510 (
            .a(out_4498),
            .b(out_4509),
            .outp(out_4510)
        );        
        

        logic [WIDTH-1:0] out_4511;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4511 (
            .in(out_4505),
            .outp(out_4511)
        );
        

        logic [WIDTH-1:0] out_4512;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4512 (
            .a(out_4501),
            .b(out_4511),
            .outp(out_4512)
        );        
        

        logic [WIDTH-1:0] out_4513;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4513 (
            .a(out_152),
            .b(out_4507),
            .outp(out_4513)
        );        
        

        logic [WIDTH-1:0] out_4514;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4514 (
            .a(out_4512),
            .b(out_4513),
            .outp(out_4514)
        );        
        

        logic [WIDTH-1:0] out_4515;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4515 (
            .a(out_4510),
            .b(out_4514),
            .outp(out_4515)
        );        
        

        logic [WIDTH-1:0] out_4516;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.7575)
        ) inst_4516 (
            .outp(out_4516)
        );
        

        logic [WIDTH-1:0] out_4517;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4517 (
            .a(out_131),
            .b(out_4516),
            .outp(out_4517)
        );        
        

        logic [WIDTH-1:0] out_4518;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4518 (
            .a(out_4517),
            .b(out_127),
            .outp(out_4518)
        );        
        

        logic [WIDTH-1:0] out_4519;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4519 (
            .a(out_4511),
            .b(out_4518),
            .outp(out_4519)
        );        
        

        logic [WIDTH-1:0] out_4520;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.195)
        ) inst_4520 (
            .outp(out_4520)
        );
        

        logic [WIDTH-1:0] out_4521;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4521 (
            .a(out_137),
            .b(out_4520),
            .outp(out_4521)
        );        
        

        logic [WIDTH-1:0] out_4522;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4522 (
            .a(out_4519),
            .b(out_4521),
            .outp(out_4522)
        );        
        

        logic [WIDTH-1:0] out_4523;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4523 (
            .a(out_4515),
            .b(out_4522),
            .outp(out_4523)
        );        
        

        logic [WIDTH-1:0] out_4524;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4524 (
            .in(out_4518),
            .outp(out_4524)
        );
        

        logic [WIDTH-1:0] out_4525;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4525 (
            .a(out_4505),
            .b(out_4524),
            .outp(out_4525)
        );        
        

        logic [WIDTH-1:0] out_4526;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4526 (
            .a(out_4520),
            .b(out_137),
            .outp(out_4526)
        );        
        

        logic [WIDTH-1:0] out_4527;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4527 (
            .a(out_4525),
            .b(out_4526),
            .outp(out_4527)
        );        
        

        logic [WIDTH-1:0] out_4528;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4528 (
            .a(out_4523),
            .b(out_4527),
            .outp(out_4528)
        );        
        

        logic [WIDTH-1:0] out_4529;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.375)
        ) inst_4529 (
            .outp(out_4529)
        );
        

        logic [WIDTH-1:0] out_4530;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4530 (
            .a(out_4529),
            .b(out_3),
            .outp(out_4530)
        );        
        

        logic [WIDTH-1:0] out_4531;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4531 (
            .in(out_4530),
            .outp(out_4531)
        );
        

        logic [WIDTH-1:0] out_4532;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.675)
        ) inst_4532 (
            .outp(out_4532)
        );
        

        logic [WIDTH-1:0] out_4533;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4533 (
            .a(out_14),
            .b(out_4532),
            .outp(out_4533)
        );        
        

        logic [WIDTH-1:0] out_4534;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4534 (
            .in(out_4533),
            .outp(out_4534)
        );
        

        logic [WIDTH-1:0] out_4535;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4535 (
            .a(out_4531),
            .b(out_4534),
            .outp(out_4535)
        );        
        

        logic [WIDTH-1:0] out_4536;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4536 (
            .in(out_4535),
            .outp(out_4536)
        );
        

        logic [WIDTH-1:0] out_4537;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4537 (
            .a(out_9),
            .b(out_4536),
            .outp(out_4537)
        );        
        

        logic [WIDTH-1:0] out_4538;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4538 (
            .a(out_4536),
            .b(out_21),
            .outp(out_4538)
        );        
        

        logic [WIDTH-1:0] out_4539;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4539 (
            .a(out_4537),
            .b(out_4538),
            .outp(out_4539)
        );        
        

        logic [WIDTH-1:0] out_4540;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4540 (
            .a(out_4528),
            .b(out_4539),
            .outp(out_4540)
        );        
        

        logic [WIDTH-1:0] out_4541;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.75)
        ) inst_4541 (
            .outp(out_4541)
        );
        

        logic [WIDTH-1:0] out_4542;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4542 (
            .a(out_4541),
            .b(out_3),
            .outp(out_4542)
        );        
        

        logic [WIDTH-1:0] out_4543;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.85)
        ) inst_4543 (
            .outp(out_4543)
        );
        

        logic [WIDTH-1:0] out_4544;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4544 (
            .a(out_4543),
            .b(out_3),
            .outp(out_4544)
        );        
        

        logic [WIDTH-1:0] out_4545;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4545 (
            .in(out_4544),
            .outp(out_4545)
        );
        

        logic [WIDTH-1:0] out_4546;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4546 (
            .a(out_4542),
            .b(out_4545),
            .outp(out_4546)
        );        
        

        logic [WIDTH-1:0] out_4547;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.725)
        ) inst_4547 (
            .outp(out_4547)
        );
        

        logic [WIDTH-1:0] out_4548;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4548 (
            .a(out_14),
            .b(out_4547),
            .outp(out_4548)
        );        
        

        logic [WIDTH-1:0] out_4549;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4549 (
            .a(out_4546),
            .b(out_4548),
            .outp(out_4549)
        );        
        

        logic [WIDTH-1:0] out_4550;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.4)
        ) inst_4550 (
            .outp(out_4550)
        );
        

        logic [WIDTH-1:0] out_4551;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4551 (
            .a(out_4550),
            .b(out_14),
            .outp(out_4551)
        );        
        

        logic [WIDTH-1:0] out_4552;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4552 (
            .a(out_4549),
            .b(out_4551),
            .outp(out_4552)
        );        
        

        logic [WIDTH-1:0] out_4553;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4553 (
            .a(out_4540),
            .b(out_4552),
            .outp(out_4553)
        );        
        

        logic [WIDTH-1:0] out_4554;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.2)
        ) inst_4554 (
            .outp(out_4554)
        );
        

        logic [WIDTH-1:0] out_4555;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4555 (
            .a(out_4554),
            .b(out_3),
            .outp(out_4555)
        );        
        

        logic [WIDTH-1:0] out_4556;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4556 (
            .a(out_3074),
            .b(out_4555),
            .outp(out_4556)
        );        
        

        logic [WIDTH-1:0] out_4557;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4557 (
            .a(out_4556),
            .b(out_4551),
            .outp(out_4557)
        );        
        

        logic [WIDTH-1:0] out_4558;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.95)
        ) inst_4558 (
            .outp(out_4558)
        );
        

        logic [WIDTH-1:0] out_4559;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4559 (
            .a(out_14),
            .b(out_4558),
            .outp(out_4559)
        );        
        

        logic [WIDTH-1:0] out_4560;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4560 (
            .a(out_4557),
            .b(out_4559),
            .outp(out_4560)
        );        
        

        logic [WIDTH-1:0] out_4561;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4561 (
            .a(out_4553),
            .b(out_4560),
            .outp(out_4561)
        );        
        

        logic [WIDTH-1:0] out_4562;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4562 (
            .a(out_3074),
            .b(out_4542),
            .outp(out_4562)
        );        
        

        logic [WIDTH-1:0] out_4563;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.025)
        ) inst_4563 (
            .outp(out_4563)
        );
        

        logic [WIDTH-1:0] out_4564;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4564 (
            .a(out_4563),
            .b(out_3),
            .outp(out_4564)
        );        
        

        logic [WIDTH-1:0] out_4565;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4565 (
            .in(out_4564),
            .outp(out_4565)
        );
        

        logic [WIDTH-1:0] out_4566;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4566 (
            .a(out_4565),
            .b(out_4534),
            .outp(out_4566)
        );        
        

        logic [WIDTH-1:0] out_4567;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4567 (
            .in(out_4566),
            .outp(out_4567)
        );
        

        logic [WIDTH-1:0] out_4568;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4568 (
            .a(out_9),
            .b(out_4567),
            .outp(out_4568)
        );        
        

        logic [WIDTH-1:0] out_4569;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4569 (
            .a(out_4562),
            .b(out_4568),
            .outp(out_4569)
        );        
        

        logic [WIDTH-1:0] out_4570;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4570 (
            .a(out_4567),
            .b(out_21),
            .outp(out_4570)
        );        
        

        logic [WIDTH-1:0] out_4571;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4571 (
            .a(out_4569),
            .b(out_4570),
            .outp(out_4571)
        );        
        

        logic [WIDTH-1:0] out_4572;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.725)
        ) inst_4572 (
            .outp(out_4572)
        );
        

        logic [WIDTH-1:0] out_4573;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4573 (
            .a(out_4572),
            .b(out_14),
            .outp(out_4573)
        );        
        

        logic [WIDTH-1:0] out_4574;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4574 (
            .a(out_4571),
            .b(out_4573),
            .outp(out_4574)
        );        
        

        logic [WIDTH-1:0] out_4575;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4575 (
            .a(out_4574),
            .b(out_4559),
            .outp(out_4575)
        );        
        

        logic [WIDTH-1:0] out_4576;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4576 (
            .a(out_4561),
            .b(out_4575),
            .outp(out_4576)
        );        
        

        logic [WIDTH-1:0] out_4577;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.825)
        ) inst_4577 (
            .outp(out_4577)
        );
        

        logic [WIDTH-1:0] out_4578;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4578 (
            .a(out_14),
            .b(out_4577),
            .outp(out_4578)
        );        
        

        logic [WIDTH-1:0] out_4579;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5)
        ) inst_4579 (
            .outp(out_4579)
        );
        

        logic [WIDTH-1:0] out_4580;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4580 (
            .a(out_4579),
            .b(out_14),
            .outp(out_4580)
        );        
        

        logic [WIDTH-1:0] out_4581;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4581 (
            .a(out_4578),
            .b(out_4580),
            .outp(out_4581)
        );        
        

        logic [WIDTH-1:0] out_4582;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.05251)
        ) inst_4582 (
            .outp(out_4582)
        );
        

        logic [WIDTH-1:0] out_4583;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4583 (
            .a(out_3),
            .b(out_4582),
            .outp(out_4583)
        );        
        

        logic [WIDTH-1:0] out_4584;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4584 (
            .a(out_4581),
            .b(out_4583),
            .outp(out_4584)
        );        
        

        logic [WIDTH-1:0] out_4585;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.95251)
        ) inst_4585 (
            .outp(out_4585)
        );
        

        logic [WIDTH-1:0] out_4586;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4586 (
            .a(out_4585),
            .b(out_3),
            .outp(out_4586)
        );        
        

        logic [WIDTH-1:0] out_4587;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4587 (
            .a(out_4584),
            .b(out_4586),
            .outp(out_4587)
        );        
        

        logic [WIDTH-1:0] out_4588;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4588 (
            .a(out_4576),
            .b(out_4587),
            .outp(out_4588)
        );        
        

        logic [WIDTH-1:0] out_4589;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.05)
        ) inst_4589 (
            .outp(out_4589)
        );
        

        logic [WIDTH-1:0] out_4590;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4590 (
            .a(out_14),
            .b(out_4589),
            .outp(out_4590)
        );        
        

        logic [WIDTH-1:0] out_4591;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4591 (
            .a(out_4580),
            .b(out_4590),
            .outp(out_4591)
        );        
        

        logic [WIDTH-1:0] out_4592;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.60251)
        ) inst_4592 (
            .outp(out_4592)
        );
        

        logic [WIDTH-1:0] out_4593;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4593 (
            .a(out_3),
            .b(out_4592),
            .outp(out_4593)
        );        
        

        logic [WIDTH-1:0] out_4594;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4594 (
            .a(out_4591),
            .b(out_4593),
            .outp(out_4594)
        );        
        

        logic [WIDTH-1:0] out_4595;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.50251)
        ) inst_4595 (
            .outp(out_4595)
        );
        

        logic [WIDTH-1:0] out_4596;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4596 (
            .a(out_4595),
            .b(out_3),
            .outp(out_4596)
        );        
        

        logic [WIDTH-1:0] out_4597;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4597 (
            .a(out_4594),
            .b(out_4596),
            .outp(out_4597)
        );        
        

        logic [WIDTH-1:0] out_4598;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4598 (
            .a(out_4588),
            .b(out_4597),
            .outp(out_4598)
        );        
        

        logic [WIDTH-1:0] out_4599;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4599 (
            .a(out_4583),
            .b(out_4590),
            .outp(out_4599)
        );        
        

        logic [WIDTH-1:0] out_4600;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4600 (
            .a(out_4599),
            .b(out_4596),
            .outp(out_4600)
        );        
        

        logic [WIDTH-1:0] out_4601;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4601 (
            .a(out_4577),
            .b(out_14),
            .outp(out_4601)
        );        
        

        logic [WIDTH-1:0] out_4602;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4602 (
            .a(out_4600),
            .b(out_4601),
            .outp(out_4602)
        );        
        

        logic [WIDTH-1:0] out_4603;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.77751)
        ) inst_4603 (
            .outp(out_4603)
        );
        

        logic [WIDTH-1:0] out_4604;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4604 (
            .a(out_3),
            .b(out_4603),
            .outp(out_4604)
        );        
        

        logic [WIDTH-1:0] out_4605;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4605 (
            .in(out_4604),
            .outp(out_4605)
        );
        

        logic [WIDTH-1:0] out_4606;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4606 (
            .a(out_4420),
            .b(out_4605),
            .outp(out_4606)
        );        
        

        logic [WIDTH-1:0] out_4607;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4607 (
            .in(out_4606),
            .outp(out_4607)
        );
        

        logic [WIDTH-1:0] out_4608;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4608 (
            .a(out_9),
            .b(out_4607),
            .outp(out_4608)
        );        
        

        logic [WIDTH-1:0] out_4609;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4609 (
            .a(out_4602),
            .b(out_4608),
            .outp(out_4609)
        );        
        

        logic [WIDTH-1:0] out_4610;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4610 (
            .a(out_4607),
            .b(out_21),
            .outp(out_4610)
        );        
        

        logic [WIDTH-1:0] out_4611;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4611 (
            .a(out_4609),
            .b(out_4610),
            .outp(out_4611)
        );        
        

        logic [WIDTH-1:0] out_4612;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4612 (
            .a(out_4598),
            .b(out_4611),
            .outp(out_4612)
        );        
        

        logic [WIDTH-1:0] out_4613;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4613 (
            .a(out_4580),
            .b(out_4419),
            .outp(out_4613)
        );        
        

        logic [WIDTH-1:0] out_4614;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1225)
        ) inst_4614 (
            .outp(out_4614)
        );
        

        logic [WIDTH-1:0] out_4615;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4615 (
            .a(out_3),
            .b(out_4614),
            .outp(out_4615)
        );        
        

        logic [WIDTH-1:0] out_4616;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4616 (
            .a(out_4613),
            .b(out_4615),
            .outp(out_4616)
        );        
        

        logic [WIDTH-1:0] out_4617;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0225)
        ) inst_4617 (
            .outp(out_4617)
        );
        

        logic [WIDTH-1:0] out_4618;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4618 (
            .a(out_4617),
            .b(out_3),
            .outp(out_4618)
        );        
        

        logic [WIDTH-1:0] out_4619;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4619 (
            .a(out_4616),
            .b(out_4618),
            .outp(out_4619)
        );        
        

        logic [WIDTH-1:0] out_4620;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4620 (
            .a(out_4612),
            .b(out_4619),
            .outp(out_4620)
        );        
        

        logic [WIDTH-1:0] out_4621;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6725)
        ) inst_4621 (
            .outp(out_4621)
        );
        

        logic [WIDTH-1:0] out_4622;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4622 (
            .a(out_3),
            .b(out_4621),
            .outp(out_4622)
        );        
        

        logic [WIDTH-1:0] out_4623;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4623 (
            .a(out_4580),
            .b(out_4622),
            .outp(out_4623)
        );        
        

        logic [WIDTH-1:0] out_4624;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5725)
        ) inst_4624 (
            .outp(out_4624)
        );
        

        logic [WIDTH-1:0] out_4625;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4625 (
            .a(out_4624),
            .b(out_3),
            .outp(out_4625)
        );        
        

        logic [WIDTH-1:0] out_4626;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4626 (
            .a(out_4623),
            .b(out_4625),
            .outp(out_4626)
        );        
        

        logic [WIDTH-1:0] out_4627;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.5)
        ) inst_4627 (
            .outp(out_4627)
        );
        

        logic [WIDTH-1:0] out_4628;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4628 (
            .a(out_14),
            .b(out_4627),
            .outp(out_4628)
        );        
        

        logic [WIDTH-1:0] out_4629;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4629 (
            .a(out_4626),
            .b(out_4628),
            .outp(out_4629)
        );        
        

        logic [WIDTH-1:0] out_4630;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4630 (
            .a(out_4620),
            .b(out_4629),
            .outp(out_4630)
        );        
        

        logic [WIDTH-1:0] out_4631;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4631 (
            .a(out_4590),
            .b(out_4625),
            .outp(out_4631)
        );        
        

        logic [WIDTH-1:0] out_4632;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8475)
        ) inst_4632 (
            .outp(out_4632)
        );
        

        logic [WIDTH-1:0] out_4633;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4633 (
            .a(out_3),
            .b(out_4632),
            .outp(out_4633)
        );        
        

        logic [WIDTH-1:0] out_4634;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4634 (
            .in(out_4633),
            .outp(out_4634)
        );
        

        logic [WIDTH-1:0] out_4635;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4635 (
            .a(out_4420),
            .b(out_4634),
            .outp(out_4635)
        );        
        

        logic [WIDTH-1:0] out_4636;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4636 (
            .in(out_4635),
            .outp(out_4636)
        );
        

        logic [WIDTH-1:0] out_4637;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4637 (
            .a(out_9),
            .b(out_4636),
            .outp(out_4637)
        );        
        

        logic [WIDTH-1:0] out_4638;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4638 (
            .a(out_4631),
            .b(out_4637),
            .outp(out_4638)
        );        
        

        logic [WIDTH-1:0] out_4639;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4639 (
            .a(out_4636),
            .b(out_21),
            .outp(out_4639)
        );        
        

        logic [WIDTH-1:0] out_4640;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4640 (
            .a(out_4638),
            .b(out_4639),
            .outp(out_4640)
        );        
        

        logic [WIDTH-1:0] out_4641;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4641 (
            .a(out_1787),
            .b(out_14),
            .outp(out_4641)
        );        
        

        logic [WIDTH-1:0] out_4642;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4642 (
            .a(out_4640),
            .b(out_4641),
            .outp(out_4642)
        );        
        

        logic [WIDTH-1:0] out_4643;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4643 (
            .a(out_4642),
            .b(out_4615),
            .outp(out_4643)
        );        
        

        logic [WIDTH-1:0] out_4644;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4644 (
            .a(out_4630),
            .b(out_4643),
            .outp(out_4644)
        );        
        

        logic [WIDTH-1:0] out_4645;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.597376)
        ) inst_4645 (
            .outp(out_4645)
        );
        

        logic [WIDTH-1:0] out_4646;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4646 (
            .a(out_4645),
            .b(out_131),
            .outp(out_4646)
        );        
        

        logic [WIDTH-1:0] out_4647;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4647 (
            .a(out_127),
            .b(out_4646),
            .outp(out_4647)
        );        
        

        logic [WIDTH-1:0] out_4648;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4648 (
            .a(out_4447),
            .b(out_4647),
            .outp(out_4648)
        );        
        

        logic [WIDTH-1:0] out_4649;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.292376)
        ) inst_4649 (
            .outp(out_4649)
        );
        

        logic [WIDTH-1:0] out_4650;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4650 (
            .a(out_4649),
            .b(out_124),
            .outp(out_4650)
        );        
        

        logic [WIDTH-1:0] out_4651;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4651 (
            .a(out_4650),
            .b(out_127),
            .outp(out_4651)
        );        
        

        logic [WIDTH-1:0] out_4652;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4652 (
            .a(out_4648),
            .b(out_4651),
            .outp(out_4652)
        );        
        

        logic [WIDTH-1:0] out_4653;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4653 (
            .a(out_4644),
            .b(out_4652),
            .outp(out_4653)
        );        
        

        logic [WIDTH-1:0] out_4654;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4654 (
            .a(out_127),
            .b(out_4650),
            .outp(out_4654)
        );        
        

        logic [WIDTH-1:0] out_4655;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4655 (
            .a(out_4460),
            .b(out_4654),
            .outp(out_4655)
        );        
        

        logic [WIDTH-1:0] out_4656;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4656 (
            .a(out_4646),
            .b(out_127),
            .outp(out_4656)
        );        
        

        logic [WIDTH-1:0] out_4657;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4657 (
            .a(out_4655),
            .b(out_4656),
            .outp(out_4657)
        );        
        

        logic [WIDTH-1:0] out_4658;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4658 (
            .a(out_4653),
            .b(out_4657),
            .outp(out_4658)
        );        
        

        logic [WIDTH-1:0] out_4659;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4659 (
            .a(out_4464),
            .b(out_4654),
            .outp(out_4659)
        );        
        

        logic [WIDTH-1:0] out_4660;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.542376)
        ) inst_4660 (
            .outp(out_4660)
        );
        

        logic [WIDTH-1:0] out_4661;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4661 (
            .a(out_4660),
            .b(out_131),
            .outp(out_4661)
        );        
        

        logic [WIDTH-1:0] out_4662;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4662 (
            .a(out_4661),
            .b(out_127),
            .outp(out_4662)
        );        
        

        logic [WIDTH-1:0] out_4663;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4663 (
            .a(out_4659),
            .b(out_4662),
            .outp(out_4663)
        );        
        

        logic [WIDTH-1:0] out_4664;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4664 (
            .a(out_4658),
            .b(out_4663),
            .outp(out_4664)
        );        
        

        logic [WIDTH-1:0] out_4665;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4665 (
            .a(out_4473),
            .b(out_4651),
            .outp(out_4665)
        );        
        

        logic [WIDTH-1:0] out_4666;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4666 (
            .a(out_127),
            .b(out_4661),
            .outp(out_4666)
        );        
        

        logic [WIDTH-1:0] out_4667;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4667 (
            .a(out_4665),
            .b(out_4666),
            .outp(out_4667)
        );        
        

        logic [WIDTH-1:0] out_4668;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4668 (
            .a(out_4664),
            .b(out_4667),
            .outp(out_4668)
        );        
        

        logic [WIDTH-1:0] out_4669;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.79238)
        ) inst_4669 (
            .outp(out_4669)
        );
        

        logic [WIDTH-1:0] out_4670;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4670 (
            .a(out_4669),
            .b(out_4477),
            .outp(out_4670)
        );        
        

        logic [WIDTH-1:0] out_4671;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4671 (
            .a(out_4447),
            .b(out_4670),
            .outp(out_4671)
        );        
        

        logic [WIDTH-1:0] out_4672;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.09738)
        ) inst_4672 (
            .outp(out_4672)
        );
        

        logic [WIDTH-1:0] out_4673;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4673 (
            .a(out_4480),
            .b(out_4672),
            .outp(out_4673)
        );        
        

        logic [WIDTH-1:0] out_4674;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4674 (
            .a(out_4671),
            .b(out_4673),
            .outp(out_4674)
        );        
        

        logic [WIDTH-1:0] out_4675;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4675 (
            .a(out_4668),
            .b(out_4674),
            .outp(out_4675)
        );        
        

        logic [WIDTH-1:0] out_4676;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4676 (
            .a(out_4672),
            .b(out_4480),
            .outp(out_4676)
        );        
        

        logic [WIDTH-1:0] out_4677;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4677 (
            .a(out_4460),
            .b(out_4676),
            .outp(out_4677)
        );        
        

        logic [WIDTH-1:0] out_4678;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4678 (
            .a(out_4477),
            .b(out_4669),
            .outp(out_4678)
        );        
        

        logic [WIDTH-1:0] out_4679;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4679 (
            .a(out_4677),
            .b(out_4678),
            .outp(out_4679)
        );        
        

        logic [WIDTH-1:0] out_4680;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4680 (
            .a(out_4675),
            .b(out_4679),
            .outp(out_4680)
        );        
        

        logic [WIDTH-1:0] out_4681;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4681 (
            .a(out_4464),
            .b(out_4676),
            .outp(out_4681)
        );        
        

        logic [WIDTH-1:0] out_4682;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.84738)
        ) inst_4682 (
            .outp(out_4682)
        );
        

        logic [WIDTH-1:0] out_4683;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4683 (
            .a(out_4477),
            .b(out_4682),
            .outp(out_4683)
        );        
        

        logic [WIDTH-1:0] out_4684;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4684 (
            .a(out_4681),
            .b(out_4683),
            .outp(out_4684)
        );        
        

        logic [WIDTH-1:0] out_4685;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4685 (
            .a(out_4680),
            .b(out_4684),
            .outp(out_4685)
        );        
        

        logic [WIDTH-1:0] out_4686;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4686 (
            .a(out_4473),
            .b(out_4673),
            .outp(out_4686)
        );        
        

        logic [WIDTH-1:0] out_4687;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4687 (
            .a(out_4682),
            .b(out_4477),
            .outp(out_4687)
        );        
        

        logic [WIDTH-1:0] out_4688;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4688 (
            .a(out_4686),
            .b(out_4687),
            .outp(out_4688)
        );        
        

        logic [WIDTH-1:0] out_4689;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4689 (
            .a(out_4685),
            .b(out_4688),
            .outp(out_4689)
        );        
        

        logic [WIDTH-1:0] out_4690;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.322376)
        ) inst_4690 (
            .outp(out_4690)
        );
        

        logic [WIDTH-1:0] out_4691;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4691 (
            .a(out_4690),
            .b(out_131),
            .outp(out_4691)
        );        
        

        logic [WIDTH-1:0] out_4692;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4692 (
            .a(out_127),
            .b(out_4691),
            .outp(out_4692)
        );        
        

        logic [WIDTH-1:0] out_4693;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4693 (
            .a(out_4447),
            .b(out_4692),
            .outp(out_4693)
        );        
        

        logic [WIDTH-1:0] out_4694;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0173756)
        ) inst_4694 (
            .outp(out_4694)
        );
        

        logic [WIDTH-1:0] out_4695;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4695 (
            .a(out_4694),
            .b(out_124),
            .outp(out_4695)
        );        
        

        logic [WIDTH-1:0] out_4696;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4696 (
            .a(out_4695),
            .b(out_127),
            .outp(out_4696)
        );        
        

        logic [WIDTH-1:0] out_4697;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4697 (
            .a(out_4693),
            .b(out_4696),
            .outp(out_4697)
        );        
        

        logic [WIDTH-1:0] out_4698;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4698 (
            .a(out_4689),
            .b(out_4697),
            .outp(out_4698)
        );        
        

        logic [WIDTH-1:0] out_4699;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4699 (
            .a(out_127),
            .b(out_4695),
            .outp(out_4699)
        );        
        

        logic [WIDTH-1:0] out_4700;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4700 (
            .a(out_4460),
            .b(out_4699),
            .outp(out_4700)
        );        
        

        logic [WIDTH-1:0] out_4701;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4701 (
            .a(out_4691),
            .b(out_127),
            .outp(out_4701)
        );        
        

        logic [WIDTH-1:0] out_4702;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4702 (
            .a(out_4700),
            .b(out_4701),
            .outp(out_4702)
        );        
        

        logic [WIDTH-1:0] out_4703;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4703 (
            .a(out_4698),
            .b(out_4702),
            .outp(out_4703)
        );        
        

        logic [WIDTH-1:0] out_4704;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4704 (
            .a(out_4464),
            .b(out_4699),
            .outp(out_4704)
        );        
        

        logic [WIDTH-1:0] out_4705;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.267376)
        ) inst_4705 (
            .outp(out_4705)
        );
        

        logic [WIDTH-1:0] out_4706;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4706 (
            .a(out_4705),
            .b(out_131),
            .outp(out_4706)
        );        
        

        logic [WIDTH-1:0] out_4707;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4707 (
            .a(out_4706),
            .b(out_127),
            .outp(out_4707)
        );        
        

        logic [WIDTH-1:0] out_4708;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4708 (
            .a(out_4704),
            .b(out_4707),
            .outp(out_4708)
        );        
        

        logic [WIDTH-1:0] out_4709;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4709 (
            .a(out_4703),
            .b(out_4708),
            .outp(out_4709)
        );        
        

        logic [WIDTH-1:0] out_4710;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4710 (
            .a(out_4473),
            .b(out_4696),
            .outp(out_4710)
        );        
        

        logic [WIDTH-1:0] out_4711;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4711 (
            .a(out_127),
            .b(out_4706),
            .outp(out_4711)
        );        
        

        logic [WIDTH-1:0] out_4712;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4712 (
            .a(out_4710),
            .b(out_4711),
            .outp(out_4712)
        );        
        

        logic [WIDTH-1:0] out_4713;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4713 (
            .a(out_4709),
            .b(out_4712),
            .outp(out_4713)
        );        
        

        logic [WIDTH-1:0] out_4714;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.51738)
        ) inst_4714 (
            .outp(out_4714)
        );
        

        logic [WIDTH-1:0] out_4715;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4715 (
            .a(out_4714),
            .b(out_4477),
            .outp(out_4715)
        );        
        

        logic [WIDTH-1:0] out_4716;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4716 (
            .a(out_4447),
            .b(out_4715),
            .outp(out_4716)
        );        
        

        logic [WIDTH-1:0] out_4717;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.82238)
        ) inst_4717 (
            .outp(out_4717)
        );
        

        logic [WIDTH-1:0] out_4718;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4718 (
            .a(out_4480),
            .b(out_4717),
            .outp(out_4718)
        );        
        

        logic [WIDTH-1:0] out_4719;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4719 (
            .a(out_4716),
            .b(out_4718),
            .outp(out_4719)
        );        
        

        logic [WIDTH-1:0] out_4720;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4720 (
            .a(out_4713),
            .b(out_4719),
            .outp(out_4720)
        );        
        

        logic [WIDTH-1:0] out_4721;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4721 (
            .a(out_4717),
            .b(out_4480),
            .outp(out_4721)
        );        
        

        logic [WIDTH-1:0] out_4722;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4722 (
            .a(out_4460),
            .b(out_4721),
            .outp(out_4722)
        );        
        

        logic [WIDTH-1:0] out_4723;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4723 (
            .a(out_4477),
            .b(out_4714),
            .outp(out_4723)
        );        
        

        logic [WIDTH-1:0] out_4724;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4724 (
            .a(out_4722),
            .b(out_4723),
            .outp(out_4724)
        );        
        

        logic [WIDTH-1:0] out_4725;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4725 (
            .a(out_4720),
            .b(out_4724),
            .outp(out_4725)
        );        
        

        logic [WIDTH-1:0] out_4726;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4726 (
            .a(out_4464),
            .b(out_4721),
            .outp(out_4726)
        );        
        

        logic [WIDTH-1:0] out_4727;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.57238)
        ) inst_4727 (
            .outp(out_4727)
        );
        

        logic [WIDTH-1:0] out_4728;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4728 (
            .a(out_4477),
            .b(out_4727),
            .outp(out_4728)
        );        
        

        logic [WIDTH-1:0] out_4729;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4729 (
            .a(out_4726),
            .b(out_4728),
            .outp(out_4729)
        );        
        

        logic [WIDTH-1:0] out_4730;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4730 (
            .a(out_4725),
            .b(out_4729),
            .outp(out_4730)
        );        
        

        logic [WIDTH-1:0] out_4731;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4731 (
            .a(out_4473),
            .b(out_4718),
            .outp(out_4731)
        );        
        

        logic [WIDTH-1:0] out_4732;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4732 (
            .a(out_4727),
            .b(out_4477),
            .outp(out_4732)
        );        
        

        logic [WIDTH-1:0] out_4733;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4733 (
            .a(out_4731),
            .b(out_4732),
            .outp(out_4733)
        );        
        

        logic [WIDTH-1:0] out_4734;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4734 (
            .a(out_4730),
            .b(out_4733),
            .outp(out_4734)
        );        
        

        logic [WIDTH-1:0] out_4735;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.0525)
        ) inst_4735 (
            .outp(out_4735)
        );
        

        logic [WIDTH-1:0] out_4736;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4736 (
            .a(out_3),
            .b(out_4735),
            .outp(out_4736)
        );        
        

        logic [WIDTH-1:0] out_4737;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4737 (
            .a(out_4409),
            .b(out_4736),
            .outp(out_4737)
        );        
        

        logic [WIDTH-1:0] out_4738;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.5525)
        ) inst_4738 (
            .outp(out_4738)
        );
        

        logic [WIDTH-1:0] out_4739;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4739 (
            .a(out_4738),
            .b(out_3),
            .outp(out_4739)
        );        
        

        logic [WIDTH-1:0] out_4740;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4740 (
            .a(out_4737),
            .b(out_4739),
            .outp(out_4740)
        );        
        

        logic [WIDTH-1:0] out_4741;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.7775)
        ) inst_4741 (
            .outp(out_4741)
        );
        

        logic [WIDTH-1:0] out_4742;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4742 (
            .a(out_3),
            .b(out_4741),
            .outp(out_4742)
        );        
        

        logic [WIDTH-1:0] out_4743;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4743 (
            .in(out_4742),
            .outp(out_4743)
        );
        

        logic [WIDTH-1:0] out_4744;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4744 (
            .a(out_4743),
            .b(out_4420),
            .outp(out_4744)
        );        
        

        logic [WIDTH-1:0] out_4745;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4745 (
            .in(out_4744),
            .outp(out_4745)
        );
        

        logic [WIDTH-1:0] out_4746;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4746 (
            .a(out_4745),
            .b(out_21),
            .outp(out_4746)
        );        
        

        logic [WIDTH-1:0] out_4747;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.30319)
        ) inst_4747 (
            .outp(out_4747)
        );
        

        logic [WIDTH-1:0] out_4748;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4748 (
            .a(out_559),
            .b(out_4747),
            .outp(out_4748)
        );        
        

        logic [WIDTH-1:0] out_4749;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4749 (
            .a(out_556),
            .b(out_4748),
            .outp(out_4749)
        );        
        

        logic [WIDTH-1:0] out_4750;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4750 (
            .a(out_4425),
            .b(out_4749),
            .outp(out_4750)
        );        
        

        logic [WIDTH-1:0] out_4751;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.92819)
        ) inst_4751 (
            .outp(out_4751)
        );
        

        logic [WIDTH-1:0] out_4752;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4752 (
            .a(out_4751),
            .b(out_2653),
            .outp(out_4752)
        );        
        

        logic [WIDTH-1:0] out_4753;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4753 (
            .a(out_4750),
            .b(out_4752),
            .outp(out_4753)
        );        
        

        logic [WIDTH-1:0] out_4754;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4754 (
            .a(out_2653),
            .b(out_4751),
            .outp(out_4754)
        );        
        

        logic [WIDTH-1:0] out_4755;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4755 (
            .a(out_4436),
            .b(out_4754),
            .outp(out_4755)
        );        
        

        logic [WIDTH-1:0] out_4756;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.30319)
        ) inst_4756 (
            .outp(out_4756)
        );
        

        logic [WIDTH-1:0] out_4757;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4757 (
            .a(out_559),
            .b(out_4756),
            .outp(out_4757)
        );        
        

        logic [WIDTH-1:0] out_4758;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4758 (
            .a(out_4757),
            .b(out_556),
            .outp(out_4758)
        );        
        

        logic [WIDTH-1:0] out_4759;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4759 (
            .a(out_4755),
            .b(out_4758),
            .outp(out_4759)
        );        
        

        logic [WIDTH-1:0] out_4760;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4760 (
            .a(out_4753),
            .b(out_4759),
            .outp(out_4760)
        );        
        

        logic [WIDTH-1:0] out_4761;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4761 (
            .in(out_4760),
            .outp(out_4761)
        );
        

        logic [WIDTH-1:0] out_4762;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4762 (
            .a(out_4746),
            .b(out_4761),
            .outp(out_4762)
        );        
        

        logic [WIDTH-1:0] out_4763;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4763 (
            .a(out_9),
            .b(out_4745),
            .outp(out_4763)
        );        
        

        logic [WIDTH-1:0] out_4764;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4764 (
            .a(out_4762),
            .b(out_4763),
            .outp(out_4764)
        );        
        

        logic [WIDTH-1:0] out_4765;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4765 (
            .a(out_4740),
            .b(out_4764),
            .outp(out_4765)
        );        
        

        logic [WIDTH-1:0] out_4766;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4766 (
            .a(out_4746),
            .b(out_4765),
            .outp(out_4766)
        );        
        

        logic [WIDTH-1:0] out_4767;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4767 (
            .a(out_4734),
            .b(out_4766),
            .outp(out_4767)
        );        
        

        logic [WIDTH-1:0] out_4768;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.6525)
        ) inst_4768 (
            .outp(out_4768)
        );
        

        logic [WIDTH-1:0] out_4769;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4769 (
            .a(out_3),
            .b(out_4768),
            .outp(out_4769)
        );        
        

        logic [WIDTH-1:0] out_4770;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4770 (
            .a(out_4613),
            .b(out_4769),
            .outp(out_4770)
        );        
        

        logic [WIDTH-1:0] out_4771;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5525)
        ) inst_4771 (
            .outp(out_4771)
        );
        

        logic [WIDTH-1:0] out_4772;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4772 (
            .a(out_4771),
            .b(out_3),
            .outp(out_4772)
        );        
        

        logic [WIDTH-1:0] out_4773;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4773 (
            .a(out_4770),
            .b(out_4772),
            .outp(out_4773)
        );        
        

        logic [WIDTH-1:0] out_4774;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4774 (
            .a(out_4767),
            .b(out_4773),
            .outp(out_4774)
        );        
        

        logic [WIDTH-1:0] out_4775;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4775 (
            .a(out_4580),
            .b(out_4628),
            .outp(out_4775)
        );        
        

        logic [WIDTH-1:0] out_4776;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.2025)
        ) inst_4776 (
            .outp(out_4776)
        );
        

        logic [WIDTH-1:0] out_4777;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4777 (
            .a(out_3),
            .b(out_4776),
            .outp(out_4777)
        );        
        

        logic [WIDTH-1:0] out_4778;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4778 (
            .a(out_4775),
            .b(out_4777),
            .outp(out_4778)
        );        
        

        logic [WIDTH-1:0] out_4779;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.1025)
        ) inst_4779 (
            .outp(out_4779)
        );
        

        logic [WIDTH-1:0] out_4780;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4780 (
            .a(out_4779),
            .b(out_3),
            .outp(out_4780)
        );        
        

        logic [WIDTH-1:0] out_4781;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4781 (
            .a(out_4778),
            .b(out_4780),
            .outp(out_4781)
        );        
        

        logic [WIDTH-1:0] out_4782;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4782 (
            .a(out_4774),
            .b(out_4781),
            .outp(out_4782)
        );        
        

        logic [WIDTH-1:0] out_4783;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4783 (
            .a(out_4590),
            .b(out_4769),
            .outp(out_4783)
        );        
        

        logic [WIDTH-1:0] out_4784;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4784 (
            .a(out_4783),
            .b(out_4780),
            .outp(out_4784)
        );        
        

        logic [WIDTH-1:0] out_4785;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4785 (
            .a(out_4784),
            .b(out_4641),
            .outp(out_4785)
        );        
        

        logic [WIDTH-1:0] out_4786;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.3775)
        ) inst_4786 (
            .outp(out_4786)
        );
        

        logic [WIDTH-1:0] out_4787;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4787 (
            .a(out_3),
            .b(out_4786),
            .outp(out_4787)
        );        
        

        logic [WIDTH-1:0] out_4788;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4788 (
            .in(out_4787),
            .outp(out_4788)
        );
        

        logic [WIDTH-1:0] out_4789;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4789 (
            .a(out_4420),
            .b(out_4788),
            .outp(out_4789)
        );        
        

        logic [WIDTH-1:0] out_4790;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4790 (
            .in(out_4789),
            .outp(out_4790)
        );
        

        logic [WIDTH-1:0] out_4791;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4791 (
            .a(out_9),
            .b(out_4790),
            .outp(out_4791)
        );        
        

        logic [WIDTH-1:0] out_4792;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4792 (
            .a(out_4785),
            .b(out_4791),
            .outp(out_4792)
        );        
        

        logic [WIDTH-1:0] out_4793;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4793 (
            .a(out_4790),
            .b(out_21),
            .outp(out_4793)
        );        
        

        logic [WIDTH-1:0] out_4794;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4794 (
            .a(out_4792),
            .b(out_4793),
            .outp(out_4794)
        );        
        

        logic [WIDTH-1:0] out_4795;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4795 (
            .a(out_4782),
            .b(out_4794),
            .outp(out_4795)
        );        
        

        logic [WIDTH-1:0] out_4796;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.300176)
        ) inst_4796 (
            .outp(out_4796)
        );
        

        logic [WIDTH-1:0] out_4797;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4797 (
            .a(out_4796),
            .b(out_1823),
            .outp(out_4797)
        );        
        

        logic [WIDTH-1:0] out_4798;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4798 (
            .a(out_4797),
            .b(out_1826),
            .outp(out_4798)
        );        
        

        logic [WIDTH-1:0] out_4799;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.26024)
        ) inst_4799 (
            .outp(out_4799)
        );
        

        logic [WIDTH-1:0] out_4800;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4800 (
            .a(out_1831),
            .b(out_4799),
            .outp(out_4800)
        );        
        

        logic [WIDTH-1:0] out_4801;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4801 (
            .a(out_4798),
            .b(out_4800),
            .outp(out_4801)
        );        
        

        logic [WIDTH-1:0] out_4802;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.80744)
        ) inst_4802 (
            .outp(out_4802)
        );
        

        logic [WIDTH-1:0] out_4803;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4803 (
            .a(out_4802),
            .b(out_1834),
            .outp(out_4803)
        );        
        

        logic [WIDTH-1:0] out_4804;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4804 (
            .a(out_4801),
            .b(out_4803),
            .outp(out_4804)
        );        
        

        logic [WIDTH-1:0] out_4805;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4805 (
            .a(out_1834),
            .b(out_4802),
            .outp(out_4805)
        );        
        

        logic [WIDTH-1:0] out_4806;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4806 (
            .a(out_4799),
            .b(out_1831),
            .outp(out_4806)
        );        
        

        logic [WIDTH-1:0] out_4807;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4807 (
            .a(out_4805),
            .b(out_4806),
            .outp(out_4807)
        );        
        

        logic [WIDTH-1:0] out_4808;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.300176)
        ) inst_4808 (
            .outp(out_4808)
        );
        

        logic [WIDTH-1:0] out_4809;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4809 (
            .a(out_4808),
            .b(out_1823),
            .outp(out_4809)
        );        
        

        logic [WIDTH-1:0] out_4810;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4810 (
            .a(out_1826),
            .b(out_4809),
            .outp(out_4810)
        );        
        

        logic [WIDTH-1:0] out_4811;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4811 (
            .a(out_4807),
            .b(out_4810),
            .outp(out_4811)
        );        
        

        logic [WIDTH-1:0] out_4812;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4812 (
            .a(out_4804),
            .b(out_4811),
            .outp(out_4812)
        );        
        

        logic [WIDTH-1:0] out_4813;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4813 (
            .in(out_4812),
            .outp(out_4813)
        );
        

        logic [WIDTH-1:0] out_4814;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.7975)
        ) inst_4814 (
            .outp(out_4814)
        );
        

        logic [WIDTH-1:0] out_4815;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4815 (
            .a(out_3),
            .b(out_4814),
            .outp(out_4815)
        );        
        

        logic [WIDTH-1:0] out_4816;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4816 (
            .in(out_4815),
            .outp(out_4816)
        );
        

        logic [WIDTH-1:0] out_4817;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4817 (
            .a(out_4420),
            .b(out_4816),
            .outp(out_4817)
        );        
        

        logic [WIDTH-1:0] out_4818;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4818 (
            .in(out_4817),
            .outp(out_4818)
        );
        

        logic [WIDTH-1:0] out_4819;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4819 (
            .a(out_9),
            .b(out_4818),
            .outp(out_4819)
        );        
        

        logic [WIDTH-1:0] out_4820;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4820 (
            .a(out_4813),
            .b(out_4819),
            .outp(out_4820)
        );        
        

        logic [WIDTH-1:0] out_4821;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4821 (
            .a(out_4818),
            .b(out_21),
            .outp(out_4821)
        );        
        

        logic [WIDTH-1:0] out_4822;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4822 (
            .a(out_4820),
            .b(out_4821),
            .outp(out_4822)
        );        
        

        logic [WIDTH-1:0] out_4823;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4823 (
            .a(out_4795),
            .b(out_4822),
            .outp(out_4823)
        );        
        

        logic [WIDTH-1:0] out_4824;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.3975)
        ) inst_4824 (
            .outp(out_4824)
        );
        

        logic [WIDTH-1:0] out_4825;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4825 (
            .a(out_3),
            .b(out_4824),
            .outp(out_4825)
        );        
        

        logic [WIDTH-1:0] out_4826;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4826 (
            .a(out_4591),
            .b(out_4825),
            .outp(out_4826)
        );        
        

        logic [WIDTH-1:0] out_4827;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2975)
        ) inst_4827 (
            .outp(out_4827)
        );
        

        logic [WIDTH-1:0] out_4828;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4828 (
            .a(out_4827),
            .b(out_3),
            .outp(out_4828)
        );        
        

        logic [WIDTH-1:0] out_4829;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4829 (
            .a(out_4826),
            .b(out_4828),
            .outp(out_4829)
        );        
        

        logic [WIDTH-1:0] out_4830;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4830 (
            .a(out_4823),
            .b(out_4829),
            .outp(out_4830)
        );        
        

        logic [WIDTH-1:0] out_4831;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2)
        ) inst_4831 (
            .outp(out_4831)
        );
        

        logic [WIDTH-1:0] out_4832;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4832 (
            .a(out_14),
            .b(out_4831),
            .outp(out_4832)
        );        
        

        logic [WIDTH-1:0] out_4833;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4833 (
            .in(out_4832),
            .outp(out_4833)
        );
        

        logic [WIDTH-1:0] out_4834;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.3475)
        ) inst_4834 (
            .outp(out_4834)
        );
        

        logic [WIDTH-1:0] out_4835;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4835 (
            .a(out_3),
            .b(out_4834),
            .outp(out_4835)
        );        
        

        logic [WIDTH-1:0] out_4836;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4836 (
            .in(out_4835),
            .outp(out_4836)
        );
        

        logic [WIDTH-1:0] out_4837;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4837 (
            .a(out_4833),
            .b(out_4836),
            .outp(out_4837)
        );        
        

        logic [WIDTH-1:0] out_4838;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4838 (
            .in(out_4837),
            .outp(out_4838)
        );
        

        logic [WIDTH-1:0] out_4839;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4839 (
            .a(out_4838),
            .b(out_460),
            .outp(out_4839)
        );        
        

        logic [WIDTH-1:0] out_4840;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4840 (
            .a(out_4830),
            .b(out_4839),
            .outp(out_4840)
        );        
        

        logic [WIDTH-1:0] out_4841;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8875)
        ) inst_4841 (
            .outp(out_4841)
        );
        

        logic [WIDTH-1:0] out_4842;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4842 (
            .a(out_14),
            .b(out_4841),
            .outp(out_4842)
        );        
        

        logic [WIDTH-1:0] out_4843;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4843 (
            .a(out_4408),
            .b(out_4842),
            .outp(out_4843)
        );        
        

        logic [WIDTH-1:0] out_4844;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5175)
        ) inst_4844 (
            .outp(out_4844)
        );
        

        logic [WIDTH-1:0] out_4845;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4845 (
            .a(out_4844),
            .b(out_260),
            .outp(out_4845)
        );        
        

        logic [WIDTH-1:0] out_4846;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4846 (
            .in(out_4845),
            .outp(out_4846)
        );
        

        logic [WIDTH-1:0] out_4847;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4847 (
            .a(out_4843),
            .b(out_4846),
            .outp(out_4847)
        );        
        

        logic [WIDTH-1:0] out_4848;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.355)
        ) inst_4848 (
            .outp(out_4848)
        );
        

        logic [WIDTH-1:0] out_4849;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4849 (
            .a(out_4848),
            .b(out_260),
            .outp(out_4849)
        );        
        

        logic [WIDTH-1:0] out_4850;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4850 (
            .a(out_4847),
            .b(out_4849),
            .outp(out_4850)
        );        
        

        logic [WIDTH-1:0] out_4851;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.885)
        ) inst_4851 (
            .outp(out_4851)
        );
        

        logic [WIDTH-1:0] out_4852;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4852 (
            .a(out_4851),
            .b(out_14),
            .outp(out_4852)
        );        
        

        logic [WIDTH-1:0] out_4853;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4853 (
            .in(out_4852),
            .outp(out_4853)
        );
        

        logic [WIDTH-1:0] out_4854;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.346667)
        ) inst_4854 (
            .outp(out_4854)
        );
        

        logic [WIDTH-1:0] out_4855;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4855 (
            .a(out_4854),
            .b(out_241),
            .outp(out_4855)
        );        
        

        logic [WIDTH-1:0] out_4856;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4856 (
            .in(out_4855),
            .outp(out_4856)
        );
        

        logic [WIDTH-1:0] out_4857;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4857 (
            .in(out_4856),
            .outp(out_4857)
        );
        

        logic [WIDTH-1:0] out_4858;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4858 (
            .a(out_4853),
            .b(out_4857),
            .outp(out_4858)
        );        
        

        logic [WIDTH-1:0] out_4859;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4859 (
            .in(out_4858),
            .outp(out_4859)
        );
        

        logic [WIDTH-1:0] out_4860;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4860 (
            .a(out_4859),
            .b(out_250),
            .outp(out_4860)
        );        
        

        logic [WIDTH-1:0] out_4861;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4861 (
            .a(out_4850),
            .b(out_4860),
            .outp(out_4861)
        );        
        

        logic [WIDTH-1:0] out_4862;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4862 (
            .in(out_4861),
            .outp(out_4862)
        );
        

        logic [WIDTH-1:0] out_4863;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4863 (
            .a(out_4841),
            .b(out_14),
            .outp(out_4863)
        );        
        

        logic [WIDTH-1:0] out_4864;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4864 (
            .in(out_4863),
            .outp(out_4864)
        );
        

        logic [WIDTH-1:0] out_4865;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4865 (
            .in(out_4846),
            .outp(out_4865)
        );
        

        logic [WIDTH-1:0] out_4866;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4866 (
            .a(out_4864),
            .b(out_4865),
            .outp(out_4866)
        );        
        

        logic [WIDTH-1:0] out_4867;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4867 (
            .in(out_4866),
            .outp(out_4867)
        );
        

        logic [WIDTH-1:0] out_4868;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4868 (
            .a(out_4867),
            .b(out_275),
            .outp(out_4868)
        );        
        

        logic [WIDTH-1:0] out_4869;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4869 (
            .a(out_4862),
            .b(out_4868),
            .outp(out_4869)
        );        
        

        logic [WIDTH-1:0] out_4870;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4870 (
            .a(out_4840),
            .b(out_4869),
            .outp(out_4870)
        );        
        

        logic [WIDTH-1:0] out_4871;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6625)
        ) inst_4871 (
            .outp(out_4871)
        );
        

        logic [WIDTH-1:0] out_4872;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4872 (
            .a(out_4871),
            .b(out_14),
            .outp(out_4872)
        );        
        

        logic [WIDTH-1:0] out_4873;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4873 (
            .a(out_4578),
            .b(out_4872),
            .outp(out_4873)
        );        
        

        logic [WIDTH-1:0] out_4874;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5175)
        ) inst_4874 (
            .outp(out_4874)
        );
        

        logic [WIDTH-1:0] out_4875;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4875 (
            .a(out_4874),
            .b(out_260),
            .outp(out_4875)
        );        
        

        logic [WIDTH-1:0] out_4876;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4876 (
            .a(out_4873),
            .b(out_4875),
            .outp(out_4876)
        );        
        

        logic [WIDTH-1:0] out_4877;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.68)
        ) inst_4877 (
            .outp(out_4877)
        );
        

        logic [WIDTH-1:0] out_4878;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4878 (
            .a(out_4877),
            .b(out_260),
            .outp(out_4878)
        );        
        

        logic [WIDTH-1:0] out_4879;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4879 (
            .in(out_4878),
            .outp(out_4879)
        );
        

        logic [WIDTH-1:0] out_4880;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4880 (
            .a(out_4876),
            .b(out_4879),
            .outp(out_4880)
        );        
        

        logic [WIDTH-1:0] out_4881;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.665)
        ) inst_4881 (
            .outp(out_4881)
        );
        

        logic [WIDTH-1:0] out_4882;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4882 (
            .a(out_14),
            .b(out_4881),
            .outp(out_4882)
        );        
        

        logic [WIDTH-1:0] out_4883;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4883 (
            .in(out_4882),
            .outp(out_4883)
        );
        

        logic [WIDTH-1:0] out_4884;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.343334)
        ) inst_4884 (
            .outp(out_4884)
        );
        

        logic [WIDTH-1:0] out_4885;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4885 (
            .a(out_4884),
            .b(out_241),
            .outp(out_4885)
        );        
        

        logic [WIDTH-1:0] out_4886;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4886 (
            .in(out_4885),
            .outp(out_4886)
        );
        

        logic [WIDTH-1:0] out_4887;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4887 (
            .a(out_4883),
            .b(out_4886),
            .outp(out_4887)
        );        
        

        logic [WIDTH-1:0] out_4888;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4888 (
            .in(out_4887),
            .outp(out_4888)
        );
        

        logic [WIDTH-1:0] out_4889;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4889 (
            .a(out_4888),
            .b(out_250),
            .outp(out_4889)
        );        
        

        logic [WIDTH-1:0] out_4890;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4890 (
            .a(out_4880),
            .b(out_4889),
            .outp(out_4890)
        );        
        

        logic [WIDTH-1:0] out_4891;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4891 (
            .in(out_4890),
            .outp(out_4891)
        );
        

        logic [WIDTH-1:0] out_4892;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4892 (
            .a(out_14),
            .b(out_4871),
            .outp(out_4892)
        );        
        

        logic [WIDTH-1:0] out_4893;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4893 (
            .in(out_4892),
            .outp(out_4893)
        );
        

        logic [WIDTH-1:0] out_4894;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4894 (
            .in(out_4875),
            .outp(out_4894)
        );
        

        logic [WIDTH-1:0] out_4895;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4895 (
            .a(out_4893),
            .b(out_4894),
            .outp(out_4895)
        );        
        

        logic [WIDTH-1:0] out_4896;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4896 (
            .in(out_4895),
            .outp(out_4896)
        );
        

        logic [WIDTH-1:0] out_4897;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4897 (
            .a(out_4896),
            .b(out_275),
            .outp(out_4897)
        );        
        

        logic [WIDTH-1:0] out_4898;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4898 (
            .a(out_4891),
            .b(out_4897),
            .outp(out_4898)
        );        
        

        logic [WIDTH-1:0] out_4899;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4899 (
            .a(out_4870),
            .b(out_4898),
            .outp(out_4899)
        );        
        

        logic [WIDTH-1:0] out_4900;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.12)
        ) inst_4900 (
            .outp(out_4900)
        );
        

        logic [WIDTH-1:0] out_4901;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4901 (
            .a(out_4900),
            .b(out_3),
            .outp(out_4901)
        );        
        

        logic [WIDTH-1:0] out_4902;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4902 (
            .a(out_4591),
            .b(out_4901),
            .outp(out_4902)
        );        
        

        logic [WIDTH-1:0] out_4903;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.22)
        ) inst_4903 (
            .outp(out_4903)
        );
        

        logic [WIDTH-1:0] out_4904;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4904 (
            .a(out_4903),
            .b(out_3),
            .outp(out_4904)
        );        
        

        logic [WIDTH-1:0] out_4905;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4905 (
            .in(out_4904),
            .outp(out_4905)
        );
        

        logic [WIDTH-1:0] out_4906;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4906 (
            .a(out_4902),
            .b(out_4905),
            .outp(out_4906)
        );        
        

        logic [WIDTH-1:0] out_4907;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4907 (
            .a(out_4899),
            .b(out_4906),
            .outp(out_4907)
        );        
        

        logic [WIDTH-1:0] out_4908;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4908 (
            .a(out_4590),
            .b(out_4641),
            .outp(out_4908)
        );        
        

        logic [WIDTH-1:0] out_4909;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.57)
        ) inst_4909 (
            .outp(out_4909)
        );
        

        logic [WIDTH-1:0] out_4910;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4910 (
            .a(out_4909),
            .b(out_3),
            .outp(out_4910)
        );        
        

        logic [WIDTH-1:0] out_4911;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4911 (
            .a(out_4908),
            .b(out_4910),
            .outp(out_4911)
        );        
        

        logic [WIDTH-1:0] out_4912;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.67)
        ) inst_4912 (
            .outp(out_4912)
        );
        

        logic [WIDTH-1:0] out_4913;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4913 (
            .a(out_4912),
            .b(out_3),
            .outp(out_4913)
        );        
        

        logic [WIDTH-1:0] out_4914;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4914 (
            .in(out_4913),
            .outp(out_4914)
        );
        

        logic [WIDTH-1:0] out_4915;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4915 (
            .a(out_4911),
            .b(out_4914),
            .outp(out_4915)
        );        
        

        logic [WIDTH-1:0] out_4916;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4916 (
            .a(out_4907),
            .b(out_4915),
            .outp(out_4916)
        );        
        

        logic [WIDTH-1:0] out_4917;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4917 (
            .a(out_4613),
            .b(out_4901),
            .outp(out_4917)
        );        
        

        logic [WIDTH-1:0] out_4918;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4918 (
            .a(out_4917),
            .b(out_4914),
            .outp(out_4918)
        );        
        

        logic [WIDTH-1:0] out_4919;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.395)
        ) inst_4919 (
            .outp(out_4919)
        );
        

        logic [WIDTH-1:0] out_4920;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4920 (
            .a(out_4919),
            .b(out_3),
            .outp(out_4920)
        );        
        

        logic [WIDTH-1:0] out_4921;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4921 (
            .in(out_4920),
            .outp(out_4921)
        );
        

        logic [WIDTH-1:0] out_4922;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4922 (
            .a(out_4420),
            .b(out_4921),
            .outp(out_4922)
        );        
        

        logic [WIDTH-1:0] out_4923;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4923 (
            .in(out_4922),
            .outp(out_4923)
        );
        

        logic [WIDTH-1:0] out_4924;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4924 (
            .a(out_9),
            .b(out_4923),
            .outp(out_4924)
        );        
        

        logic [WIDTH-1:0] out_4925;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4925 (
            .a(out_4918),
            .b(out_4924),
            .outp(out_4925)
        );        
        

        logic [WIDTH-1:0] out_4926;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4926 (
            .a(out_4923),
            .b(out_21),
            .outp(out_4926)
        );        
        

        logic [WIDTH-1:0] out_4927;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4927 (
            .a(out_4925),
            .b(out_4926),
            .outp(out_4927)
        );        
        

        logic [WIDTH-1:0] out_4928;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4928 (
            .a(out_4916),
            .b(out_4927),
            .outp(out_4928)
        );        
        

        logic [WIDTH-1:0] out_4929;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.85)
        ) inst_4929 (
            .outp(out_4929)
        );
        

        logic [WIDTH-1:0] out_4930;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4930 (
            .a(out_14),
            .b(out_4929),
            .outp(out_4930)
        );        
        

        logic [WIDTH-1:0] out_4931;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4931 (
            .a(out_4580),
            .b(out_4930),
            .outp(out_4931)
        );        
        

        logic [WIDTH-1:0] out_4932;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.77)
        ) inst_4932 (
            .outp(out_4932)
        );
        

        logic [WIDTH-1:0] out_4933;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4933 (
            .a(out_4932),
            .b(out_3),
            .outp(out_4933)
        );        
        

        logic [WIDTH-1:0] out_4934;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4934 (
            .a(out_4931),
            .b(out_4933),
            .outp(out_4934)
        );        
        

        logic [WIDTH-1:0] out_4935;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.87)
        ) inst_4935 (
            .outp(out_4935)
        );
        

        logic [WIDTH-1:0] out_4936;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4936 (
            .a(out_4935),
            .b(out_3),
            .outp(out_4936)
        );        
        

        logic [WIDTH-1:0] out_4937;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4937 (
            .in(out_4936),
            .outp(out_4937)
        );
        

        logic [WIDTH-1:0] out_4938;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4938 (
            .a(out_4934),
            .b(out_4937),
            .outp(out_4938)
        );        
        

        logic [WIDTH-1:0] out_4939;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4939 (
            .a(out_4928),
            .b(out_4938),
            .outp(out_4939)
        );        
        

        logic [WIDTH-1:0] out_4940;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.02)
        ) inst_4940 (
            .outp(out_4940)
        );
        

        logic [WIDTH-1:0] out_4941;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4941 (
            .a(out_4940),
            .b(out_3),
            .outp(out_4941)
        );        
        

        logic [WIDTH-1:0] out_4942;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4942 (
            .a(out_4931),
            .b(out_4941),
            .outp(out_4942)
        );        
        

        logic [WIDTH-1:0] out_4943;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4943 (
            .a(out_926),
            .b(out_3),
            .outp(out_4943)
        );        
        

        logic [WIDTH-1:0] out_4944;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4944 (
            .in(out_4943),
            .outp(out_4944)
        );
        

        logic [WIDTH-1:0] out_4945;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4945 (
            .a(out_4942),
            .b(out_4944),
            .outp(out_4945)
        );        
        

        logic [WIDTH-1:0] out_4946;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4946 (
            .a(out_4939),
            .b(out_4945),
            .outp(out_4946)
        );        
        

        logic [WIDTH-1:0] out_4947;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0958748)
        ) inst_4947 (
            .outp(out_4947)
        );
        

        logic [WIDTH-1:0] out_4948;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4948 (
            .a(out_4947),
            .b(out_1891),
            .outp(out_4948)
        );        
        

        logic [WIDTH-1:0] out_4949;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4949 (
            .a(out_4948),
            .b(out_137),
            .outp(out_4949)
        );        
        

        logic [WIDTH-1:0] out_4950;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.26444)
        ) inst_4950 (
            .outp(out_4950)
        );
        

        logic [WIDTH-1:0] out_4951;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4951 (
            .a(out_4950),
            .b(out_4052),
            .outp(out_4951)
        );        
        

        logic [WIDTH-1:0] out_4952;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4952 (
            .a(out_4949),
            .b(out_4951),
            .outp(out_4952)
        );        
        

        logic [WIDTH-1:0] out_4953;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.55781)
        ) inst_4953 (
            .outp(out_4953)
        );
        

        logic [WIDTH-1:0] out_4954;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4954 (
            .a(out_1907),
            .b(out_4953),
            .outp(out_4954)
        );        
        

        logic [WIDTH-1:0] out_4955;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4955 (
            .a(out_1904),
            .b(out_4954),
            .outp(out_4955)
        );        
        

        logic [WIDTH-1:0] out_4956;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4956 (
            .a(out_4952),
            .b(out_4955),
            .outp(out_4956)
        );        
        

        logic [WIDTH-1:0] out_4957;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4957 (
            .a(out_4954),
            .b(out_1904),
            .outp(out_4957)
        );        
        

        logic [WIDTH-1:0] out_4958;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.26444)
        ) inst_4958 (
            .outp(out_4958)
        );
        

        logic [WIDTH-1:0] out_4959;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4959 (
            .a(out_4052),
            .b(out_4958),
            .outp(out_4959)
        );        
        

        logic [WIDTH-1:0] out_4960;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4960 (
            .a(out_4957),
            .b(out_4959),
            .outp(out_4960)
        );        
        

        logic [WIDTH-1:0] out_4961;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.095875)
        ) inst_4961 (
            .outp(out_4961)
        );
        

        logic [WIDTH-1:0] out_4962;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4962 (
            .a(out_4961),
            .b(out_1891),
            .outp(out_4962)
        );        
        

        logic [WIDTH-1:0] out_4963;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4963 (
            .a(out_137),
            .b(out_4962),
            .outp(out_4963)
        );        
        

        logic [WIDTH-1:0] out_4964;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4964 (
            .a(out_4960),
            .b(out_4963),
            .outp(out_4964)
        );        
        

        logic [WIDTH-1:0] out_4965;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4965 (
            .a(out_4956),
            .b(out_4964),
            .outp(out_4965)
        );        
        

        logic [WIDTH-1:0] out_4966;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4966 (
            .in(out_4965),
            .outp(out_4966)
        );
        

        logic [WIDTH-1:0] out_4967;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.575)
        ) inst_4967 (
            .outp(out_4967)
        );
        

        logic [WIDTH-1:0] out_4968;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4968 (
            .a(out_14),
            .b(out_4967),
            .outp(out_4968)
        );        
        

        logic [WIDTH-1:0] out_4969;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4969 (
            .a(out_4966),
            .b(out_4968),
            .outp(out_4969)
        );        
        

        logic [WIDTH-1:0] out_4970;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.35)
        ) inst_4970 (
            .outp(out_4970)
        );
        

        logic [WIDTH-1:0] out_4971;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4971 (
            .a(out_4970),
            .b(out_14),
            .outp(out_4971)
        );        
        

        logic [WIDTH-1:0] out_4972;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4972 (
            .a(out_4969),
            .b(out_4971),
            .outp(out_4972)
        );        
        

        logic [WIDTH-1:0] out_4973;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5475)
        ) inst_4973 (
            .outp(out_4973)
        );
        

        logic [WIDTH-1:0] out_4974;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4974 (
            .a(out_3),
            .b(out_4973),
            .outp(out_4974)
        );        
        

        logic [WIDTH-1:0] out_4975;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4975 (
            .a(out_4972),
            .b(out_4974),
            .outp(out_4975)
        );        
        

        logic [WIDTH-1:0] out_4976;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.3975)
        ) inst_4976 (
            .outp(out_4976)
        );
        

        logic [WIDTH-1:0] out_4977;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4977 (
            .a(out_4976),
            .b(out_3),
            .outp(out_4977)
        );        
        

        logic [WIDTH-1:0] out_4978;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4978 (
            .a(out_4975),
            .b(out_4977),
            .outp(out_4978)
        );        
        

        logic [WIDTH-1:0] out_4979;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.858333)
        ) inst_4979 (
            .outp(out_4979)
        );
        

        logic [WIDTH-1:0] out_4980;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4980 (
            .a(out_1933),
            .b(out_4979),
            .outp(out_4980)
        );        
        

        logic [WIDTH-1:0] out_4981;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4981 (
            .in(out_4980),
            .outp(out_4981)
        );
        

        logic [WIDTH-1:0] out_4982;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4725)
        ) inst_4982 (
            .outp(out_4982)
        );
        

        logic [WIDTH-1:0] out_4983;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4983 (
            .a(out_3),
            .b(out_4982),
            .outp(out_4983)
        );        
        

        logic [WIDTH-1:0] out_4984;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4984 (
            .in(out_4983),
            .outp(out_4984)
        );
        

        logic [WIDTH-1:0] out_4985;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4985 (
            .a(out_4981),
            .b(out_4984),
            .outp(out_4985)
        );        
        

        logic [WIDTH-1:0] out_4986;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4986 (
            .in(out_4985),
            .outp(out_4986)
        );
        

        logic [WIDTH-1:0] out_4987;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4987 (
            .a(out_4986),
            .b(out_460),
            .outp(out_4987)
        );        
        

        logic [WIDTH-1:0] out_4988;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4988 (
            .a(out_4978),
            .b(out_4987),
            .outp(out_4988)
        );        
        

        logic [WIDTH-1:0] out_4989;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4989 (
            .a(out_4946),
            .b(out_4988),
            .outp(out_4989)
        );        
        

        logic [WIDTH-1:0] out_4990;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4990 (
            .in(out_4968),
            .outp(out_4990)
        );
        

        logic [WIDTH-1:0] out_4991;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4975)
        ) inst_4991 (
            .outp(out_4991)
        );
        

        logic [WIDTH-1:0] out_4992;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4992 (
            .a(out_3),
            .b(out_4991),
            .outp(out_4992)
        );        
        

        logic [WIDTH-1:0] out_4993;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4993 (
            .in(out_4992),
            .outp(out_4993)
        );
        

        logic [WIDTH-1:0] out_4994;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4994 (
            .a(out_4990),
            .b(out_4993),
            .outp(out_4994)
        );        
        

        logic [WIDTH-1:0] out_4995;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4995 (
            .in(out_4994),
            .outp(out_4995)
        );
        

        logic [WIDTH-1:0] out_4996;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4996 (
            .a(out_4995),
            .b(out_460),
            .outp(out_4996)
        );        
        

        logic [WIDTH-1:0] out_4997;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4997 (
            .a(out_4989),
            .b(out_4996),
            .outp(out_4997)
        );        
        

        logic [WIDTH-1:0] out_4998;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.737225)
        ) inst_4998 (
            .outp(out_4998)
        );
        

        logic [WIDTH-1:0] out_4999;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_4999 (
            .a(out_4998),
            .b(out_1826),
            .outp(out_4999)
        );        
        

        logic [WIDTH-1:0] out_5000;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5000 (
            .a(out_1823),
            .b(out_4999),
            .outp(out_5000)
        );        
        

        logic [WIDTH-1:0] out_5001;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.203962)
        ) inst_5001 (
            .outp(out_5001)
        );
        

        logic [WIDTH-1:0] out_5002;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5002 (
            .a(out_1831),
            .b(out_5001),
            .outp(out_5002)
        );        
        

        logic [WIDTH-1:0] out_5003;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5003 (
            .a(out_5000),
            .b(out_5002),
            .outp(out_5003)
        );        
        

        logic [WIDTH-1:0] out_5004;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.788562)
        ) inst_5004 (
            .outp(out_5004)
        );
        

        logic [WIDTH-1:0] out_5005;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5005 (
            .a(out_5004),
            .b(out_1834),
            .outp(out_5005)
        );        
        

        logic [WIDTH-1:0] out_5006;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5006 (
            .a(out_5003),
            .b(out_5005),
            .outp(out_5006)
        );        
        

        logic [WIDTH-1:0] out_5007;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5007 (
            .a(out_1834),
            .b(out_5004),
            .outp(out_5007)
        );        
        

        logic [WIDTH-1:0] out_5008;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5008 (
            .a(out_5001),
            .b(out_1831),
            .outp(out_5008)
        );        
        

        logic [WIDTH-1:0] out_5009;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5009 (
            .a(out_5007),
            .b(out_5008),
            .outp(out_5009)
        );        
        

        logic [WIDTH-1:0] out_5010;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.737225)
        ) inst_5010 (
            .outp(out_5010)
        );
        

        logic [WIDTH-1:0] out_5011;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5011 (
            .a(out_5010),
            .b(out_1826),
            .outp(out_5011)
        );        
        

        logic [WIDTH-1:0] out_5012;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5012 (
            .a(out_5011),
            .b(out_1823),
            .outp(out_5012)
        );        
        

        logic [WIDTH-1:0] out_5013;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5013 (
            .a(out_5009),
            .b(out_5012),
            .outp(out_5013)
        );        
        

        logic [WIDTH-1:0] out_5014;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5014 (
            .a(out_5006),
            .b(out_5013),
            .outp(out_5014)
        );        
        

        logic [WIDTH-1:0] out_5015;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5015 (
            .in(out_5014),
            .outp(out_5015)
        );
        

        logic [WIDTH-1:0] out_5016;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0924997)
        ) inst_5016 (
            .outp(out_5016)
        );
        

        logic [WIDTH-1:0] out_5017;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5017 (
            .a(out_3),
            .b(out_5016),
            .outp(out_5017)
        );        
        

        logic [WIDTH-1:0] out_5018;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5018 (
            .in(out_5017),
            .outp(out_5018)
        );
        

        logic [WIDTH-1:0] out_5019;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5019 (
            .a(out_4420),
            .b(out_5018),
            .outp(out_5019)
        );        
        

        logic [WIDTH-1:0] out_5020;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5020 (
            .in(out_5019),
            .outp(out_5020)
        );
        

        logic [WIDTH-1:0] out_5021;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5021 (
            .a(out_9),
            .b(out_5020),
            .outp(out_5021)
        );        
        

        logic [WIDTH-1:0] out_5022;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5022 (
            .a(out_5015),
            .b(out_5021),
            .outp(out_5022)
        );        
        

        logic [WIDTH-1:0] out_5023;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5023 (
            .a(out_5020),
            .b(out_21),
            .outp(out_5023)
        );        
        

        logic [WIDTH-1:0] out_5024;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5024 (
            .a(out_5022),
            .b(out_5023),
            .outp(out_5024)
        );        
        

        logic [WIDTH-1:0] out_5025;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5025 (
            .a(out_4997),
            .b(out_5024),
            .outp(out_5025)
        );        
        

        logic [WIDTH-1:0] out_5026;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.3075)
        ) inst_5026 (
            .outp(out_5026)
        );
        

        logic [WIDTH-1:0] out_5027;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5027 (
            .a(out_5026),
            .b(out_3),
            .outp(out_5027)
        );        
        

        logic [WIDTH-1:0] out_5028;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5028 (
            .a(out_4591),
            .b(out_5027),
            .outp(out_5028)
        );        
        

        logic [WIDTH-1:0] out_5029;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4075)
        ) inst_5029 (
            .outp(out_5029)
        );
        

        logic [WIDTH-1:0] out_5030;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5030 (
            .a(out_5029),
            .b(out_3),
            .outp(out_5030)
        );        
        

        logic [WIDTH-1:0] out_5031;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5031 (
            .in(out_5030),
            .outp(out_5031)
        );
        

        logic [WIDTH-1:0] out_5032;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5032 (
            .a(out_5028),
            .b(out_5031),
            .outp(out_5032)
        );        
        

        logic [WIDTH-1:0] out_5033;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5033 (
            .a(out_5025),
            .b(out_5032),
            .outp(out_5033)
        );        
        

        logic [WIDTH-1:0] out_5034;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.357501)
        ) inst_5034 (
            .outp(out_5034)
        );
        

        logic [WIDTH-1:0] out_5035;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5035 (
            .a(out_5034),
            .b(out_3),
            .outp(out_5035)
        );        
        

        logic [WIDTH-1:0] out_5036;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5036 (
            .in(out_5035),
            .outp(out_5036)
        );
        

        logic [WIDTH-1:0] out_5037;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5037 (
            .a(out_4833),
            .b(out_5036),
            .outp(out_5037)
        );        
        

        logic [WIDTH-1:0] out_5038;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5038 (
            .in(out_5037),
            .outp(out_5038)
        );
        

        logic [WIDTH-1:0] out_5039;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5039 (
            .a(out_5038),
            .b(out_460),
            .outp(out_5039)
        );        
        

        logic [WIDTH-1:0] out_5040;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5040 (
            .a(out_5033),
            .b(out_5039),
            .outp(out_5040)
        );        
        

        logic [WIDTH-1:0] out_5041;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.845)
        ) inst_5041 (
            .outp(out_5041)
        );
        

        logic [WIDTH-1:0] out_5042;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5042 (
            .a(out_5041),
            .b(out_3),
            .outp(out_5042)
        );        
        

        logic [WIDTH-1:0] out_5043;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5043 (
            .a(out_4775),
            .b(out_5042),
            .outp(out_5043)
        );        
        

        logic [WIDTH-1:0] out_5044;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.945)
        ) inst_5044 (
            .outp(out_5044)
        );
        

        logic [WIDTH-1:0] out_5045;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5045 (
            .a(out_5044),
            .b(out_3),
            .outp(out_5045)
        );        
        

        logic [WIDTH-1:0] out_5046;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5046 (
            .in(out_5045),
            .outp(out_5046)
        );
        

        logic [WIDTH-1:0] out_5047;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5047 (
            .a(out_5043),
            .b(out_5046),
            .outp(out_5047)
        );        
        

        logic [WIDTH-1:0] out_5048;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5048 (
            .a(out_5040),
            .b(out_5047),
            .outp(out_5048)
        );        
        

        logic [WIDTH-1:0] out_5049;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.07)
        ) inst_5049 (
            .outp(out_5049)
        );
        

        logic [WIDTH-1:0] out_5050;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5050 (
            .a(out_5049),
            .b(out_3),
            .outp(out_5050)
        );        
        

        logic [WIDTH-1:0] out_5051;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5051 (
            .a(out_4581),
            .b(out_5050),
            .outp(out_5051)
        );        
        

        logic [WIDTH-1:0] out_5052;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.17)
        ) inst_5052 (
            .outp(out_5052)
        );
        

        logic [WIDTH-1:0] out_5053;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5053 (
            .a(out_5052),
            .b(out_3),
            .outp(out_5053)
        );        
        

        logic [WIDTH-1:0] out_5054;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5054 (
            .in(out_5053),
            .outp(out_5054)
        );
        

        logic [WIDTH-1:0] out_5055;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5055 (
            .a(out_5051),
            .b(out_5054),
            .outp(out_5055)
        );        
        

        logic [WIDTH-1:0] out_5056;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5056 (
            .a(out_5048),
            .b(out_5055),
            .outp(out_5056)
        );        
        

        logic [WIDTH-1:0] out_5057;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.52)
        ) inst_5057 (
            .outp(out_5057)
        );
        

        logic [WIDTH-1:0] out_5058;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5058 (
            .a(out_5057),
            .b(out_3),
            .outp(out_5058)
        );        
        

        logic [WIDTH-1:0] out_5059;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5059 (
            .a(out_4591),
            .b(out_5058),
            .outp(out_5059)
        );        
        

        logic [WIDTH-1:0] out_5060;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.62)
        ) inst_5060 (
            .outp(out_5060)
        );
        

        logic [WIDTH-1:0] out_5061;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5061 (
            .a(out_5060),
            .b(out_3),
            .outp(out_5061)
        );        
        

        logic [WIDTH-1:0] out_5062;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5062 (
            .in(out_5061),
            .outp(out_5062)
        );
        

        logic [WIDTH-1:0] out_5063;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5063 (
            .a(out_5059),
            .b(out_5062),
            .outp(out_5063)
        );        
        

        logic [WIDTH-1:0] out_5064;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5064 (
            .a(out_5056),
            .b(out_5063),
            .outp(out_5064)
        );        
        

        logic [WIDTH-1:0] out_5065;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5065 (
            .a(out_4590),
            .b(out_4601),
            .outp(out_5065)
        );        
        

        logic [WIDTH-1:0] out_5066;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5066 (
            .a(out_5065),
            .b(out_5050),
            .outp(out_5066)
        );        
        

        logic [WIDTH-1:0] out_5067;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5067 (
            .a(out_5066),
            .b(out_5062),
            .outp(out_5067)
        );        
        

        logic [WIDTH-1:0] out_5068;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.345)
        ) inst_5068 (
            .outp(out_5068)
        );
        

        logic [WIDTH-1:0] out_5069;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5069 (
            .a(out_5068),
            .b(out_3),
            .outp(out_5069)
        );        
        

        logic [WIDTH-1:0] out_5070;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5070 (
            .in(out_5069),
            .outp(out_5070)
        );
        

        logic [WIDTH-1:0] out_5071;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5071 (
            .a(out_4420),
            .b(out_5070),
            .outp(out_5071)
        );        
        

        logic [WIDTH-1:0] out_5072;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5072 (
            .in(out_5071),
            .outp(out_5072)
        );
        

        logic [WIDTH-1:0] out_5073;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5073 (
            .a(out_9),
            .b(out_5072),
            .outp(out_5073)
        );        
        

        logic [WIDTH-1:0] out_5074;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5074 (
            .a(out_5067),
            .b(out_5073),
            .outp(out_5074)
        );        
        

        logic [WIDTH-1:0] out_5075;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5075 (
            .a(out_5072),
            .b(out_21),
            .outp(out_5075)
        );        
        

        logic [WIDTH-1:0] out_5076;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5076 (
            .a(out_5074),
            .b(out_5075),
            .outp(out_5076)
        );        
        

        logic [WIDTH-1:0] out_5077;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5077 (
            .a(out_5064),
            .b(out_5076),
            .outp(out_5077)
        );        
        

        logic [WIDTH-1:0] out_5078;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.72)
        ) inst_5078 (
            .outp(out_5078)
        );
        

        logic [WIDTH-1:0] out_5079;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5079 (
            .a(out_5078),
            .b(out_3),
            .outp(out_5079)
        );        
        

        logic [WIDTH-1:0] out_5080;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5080 (
            .a(out_4409),
            .b(out_5079),
            .outp(out_5080)
        );        
        

        logic [WIDTH-1:0] out_5081;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.22)
        ) inst_5081 (
            .outp(out_5081)
        );
        

        logic [WIDTH-1:0] out_5082;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5082 (
            .a(out_5081),
            .b(out_3),
            .outp(out_5082)
        );        
        

        logic [WIDTH-1:0] out_5083;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5083 (
            .in(out_5082),
            .outp(out_5083)
        );
        

        logic [WIDTH-1:0] out_5084;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5084 (
            .a(out_5080),
            .b(out_5083),
            .outp(out_5084)
        );        
        

        logic [WIDTH-1:0] out_5085;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.995)
        ) inst_5085 (
            .outp(out_5085)
        );
        

        logic [WIDTH-1:0] out_5086;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5086 (
            .a(out_5085),
            .b(out_3),
            .outp(out_5086)
        );        
        

        logic [WIDTH-1:0] out_5087;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5087 (
            .in(out_5086),
            .outp(out_5087)
        );
        

        logic [WIDTH-1:0] out_5088;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5088 (
            .a(out_4420),
            .b(out_5087),
            .outp(out_5088)
        );        
        

        logic [WIDTH-1:0] out_5089;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5089 (
            .in(out_5088),
            .outp(out_5089)
        );
        

        logic [WIDTH-1:0] out_5090;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5090 (
            .a(out_5089),
            .b(out_21),
            .outp(out_5090)
        );        
        

        logic [WIDTH-1:0] out_5091;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.65925)
        ) inst_5091 (
            .outp(out_5091)
        );
        

        logic [WIDTH-1:0] out_5092;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5092 (
            .a(out_5091),
            .b(out_556),
            .outp(out_5092)
        );        
        

        logic [WIDTH-1:0] out_5093;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5093 (
            .a(out_5092),
            .b(out_559),
            .outp(out_5093)
        );        
        

        logic [WIDTH-1:0] out_5094;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5094 (
            .a(out_4425),
            .b(out_5093),
            .outp(out_5094)
        );        
        

        logic [WIDTH-1:0] out_5095;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.03425)
        ) inst_5095 (
            .outp(out_5095)
        );
        

        logic [WIDTH-1:0] out_5096;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5096 (
            .a(out_5095),
            .b(out_556),
            .outp(out_5096)
        );        
        

        logic [WIDTH-1:0] out_5097;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5097 (
            .a(out_5096),
            .b(out_566),
            .outp(out_5097)
        );        
        

        logic [WIDTH-1:0] out_5098;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5098 (
            .in(out_5097),
            .outp(out_5098)
        );
        

        logic [WIDTH-1:0] out_5099;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5099 (
            .a(out_5094),
            .b(out_5098),
            .outp(out_5099)
        );        
        

        logic [WIDTH-1:0] out_5100;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5100 (
            .a(out_4436),
            .b(out_5097),
            .outp(out_5100)
        );        
        

        logic [WIDTH-1:0] out_5101;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5101 (
            .a(out_559),
            .b(out_5092),
            .outp(out_5101)
        );        
        

        logic [WIDTH-1:0] out_5102;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5102 (
            .a(out_5100),
            .b(out_5101),
            .outp(out_5102)
        );        
        

        logic [WIDTH-1:0] out_5103;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5103 (
            .a(out_5099),
            .b(out_5102),
            .outp(out_5103)
        );        
        

        logic [WIDTH-1:0] out_5104;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5104 (
            .in(out_5103),
            .outp(out_5104)
        );
        

        logic [WIDTH-1:0] out_5105;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5105 (
            .a(out_5090),
            .b(out_5104),
            .outp(out_5105)
        );        
        

        logic [WIDTH-1:0] out_5106;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5106 (
            .a(out_9),
            .b(out_5089),
            .outp(out_5106)
        );        
        

        logic [WIDTH-1:0] out_5107;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5107 (
            .a(out_5105),
            .b(out_5106),
            .outp(out_5107)
        );        
        

        logic [WIDTH-1:0] out_5108;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5108 (
            .a(out_5084),
            .b(out_5107),
            .outp(out_5108)
        );        
        

        logic [WIDTH-1:0] out_5109;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5109 (
            .a(out_5090),
            .b(out_5108),
            .outp(out_5109)
        );        
        

        logic [WIDTH-1:0] out_5110;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5110 (
            .a(out_5077),
            .b(out_5109),
            .outp(out_5110)
        );        
        

        logic [WIDTH-1:0] out_5111;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.716)
        ) inst_5111 (
            .outp(out_5111)
        );
        

        logic [WIDTH-1:0] out_5112;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5112 (
            .a(out_5111),
            .b(out_127),
            .outp(out_5112)
        );        
        

        logic [WIDTH-1:0] out_5113;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5113 (
            .a(out_5112),
            .b(out_131),
            .outp(out_5113)
        );        
        

        logic [WIDTH-1:0] out_5114;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5114 (
            .a(out_4447),
            .b(out_5113),
            .outp(out_5114)
        );        
        

        logic [WIDTH-1:0] out_5115;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.021)
        ) inst_5115 (
            .outp(out_5115)
        );
        

        logic [WIDTH-1:0] out_5116;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5116 (
            .a(out_5115),
            .b(out_127),
            .outp(out_5116)
        );        
        

        logic [WIDTH-1:0] out_5117;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5117 (
            .a(out_124),
            .b(out_5116),
            .outp(out_5117)
        );        
        

        logic [WIDTH-1:0] out_5118;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5118 (
            .a(out_5114),
            .b(out_5117),
            .outp(out_5118)
        );        
        

        logic [WIDTH-1:0] out_5119;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5119 (
            .a(out_5110),
            .b(out_5118),
            .outp(out_5119)
        );        
        

        logic [WIDTH-1:0] out_5120;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5120 (
            .a(out_5116),
            .b(out_124),
            .outp(out_5120)
        );        
        

        logic [WIDTH-1:0] out_5121;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5121 (
            .a(out_4460),
            .b(out_5120),
            .outp(out_5121)
        );        
        

        logic [WIDTH-1:0] out_5122;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5122 (
            .a(out_131),
            .b(out_5112),
            .outp(out_5122)
        );        
        

        logic [WIDTH-1:0] out_5123;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5123 (
            .a(out_5121),
            .b(out_5122),
            .outp(out_5123)
        );        
        

        logic [WIDTH-1:0] out_5124;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5124 (
            .a(out_5119),
            .b(out_5123),
            .outp(out_5124)
        );        
        

        logic [WIDTH-1:0] out_5125;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5125 (
            .a(out_4464),
            .b(out_5120),
            .outp(out_5125)
        );        
        

        logic [WIDTH-1:0] out_5126;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.771)
        ) inst_5126 (
            .outp(out_5126)
        );
        

        logic [WIDTH-1:0] out_5127;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5127 (
            .a(out_5126),
            .b(out_127),
            .outp(out_5127)
        );        
        

        logic [WIDTH-1:0] out_5128;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5128 (
            .a(out_131),
            .b(out_5127),
            .outp(out_5128)
        );        
        

        logic [WIDTH-1:0] out_5129;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5129 (
            .a(out_5125),
            .b(out_5128),
            .outp(out_5129)
        );        
        

        logic [WIDTH-1:0] out_5130;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5130 (
            .a(out_5124),
            .b(out_5129),
            .outp(out_5130)
        );        
        

        logic [WIDTH-1:0] out_5131;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5131 (
            .a(out_4473),
            .b(out_5117),
            .outp(out_5131)
        );        
        

        logic [WIDTH-1:0] out_5132;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5132 (
            .a(out_5127),
            .b(out_131),
            .outp(out_5132)
        );        
        

        logic [WIDTH-1:0] out_5133;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5133 (
            .a(out_5131),
            .b(out_5132),
            .outp(out_5133)
        );        
        

        logic [WIDTH-1:0] out_5134;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5134 (
            .a(out_5130),
            .b(out_5133),
            .outp(out_5134)
        );        
        

        logic [WIDTH-1:0] out_5135;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.521)
        ) inst_5135 (
            .outp(out_5135)
        );
        

        logic [WIDTH-1:0] out_5136;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5136 (
            .a(out_131),
            .b(out_5135),
            .outp(out_5136)
        );        
        

        logic [WIDTH-1:0] out_5137;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5137 (
            .a(out_5136),
            .b(out_127),
            .outp(out_5137)
        );        
        

        logic [WIDTH-1:0] out_5138;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5138 (
            .in(out_5137),
            .outp(out_5138)
        );
        

        logic [WIDTH-1:0] out_5139;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5139 (
            .a(out_4447),
            .b(out_5138),
            .outp(out_5139)
        );        
        

        logic [WIDTH-1:0] out_5140;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.216)
        ) inst_5140 (
            .outp(out_5140)
        );
        

        logic [WIDTH-1:0] out_5141;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5141 (
            .a(out_5140),
            .b(out_124),
            .outp(out_5141)
        );        
        

        logic [WIDTH-1:0] out_5142;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5142 (
            .a(out_5141),
            .b(out_127),
            .outp(out_5142)
        );        
        

        logic [WIDTH-1:0] out_5143;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5143 (
            .a(out_5139),
            .b(out_5142),
            .outp(out_5143)
        );        
        

        logic [WIDTH-1:0] out_5144;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5144 (
            .a(out_5134),
            .b(out_5143),
            .outp(out_5144)
        );        
        

        logic [WIDTH-1:0] out_5145;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.025)
        ) inst_5145 (
            .outp(out_5145)
        );
        

        logic [WIDTH-1:0] out_5146;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5146 (
            .a(out_14),
            .b(out_5145),
            .outp(out_5146)
        );        
        

        logic [WIDTH-1:0] out_5147;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5147 (
            .a(out_4580),
            .b(out_5146),
            .outp(out_5147)
        );        
        

        logic [WIDTH-1:0] out_5148;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.27)
        ) inst_5148 (
            .outp(out_5148)
        );
        

        logic [WIDTH-1:0] out_5149;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5149 (
            .a(out_5148),
            .b(out_3),
            .outp(out_5149)
        );        
        

        logic [WIDTH-1:0] out_5150;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5150 (
            .a(out_5147),
            .b(out_5149),
            .outp(out_5150)
        );        
        

        logic [WIDTH-1:0] out_5151;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.37)
        ) inst_5151 (
            .outp(out_5151)
        );
        

        logic [WIDTH-1:0] out_5152;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5152 (
            .a(out_5151),
            .b(out_3),
            .outp(out_5152)
        );        
        

        logic [WIDTH-1:0] out_5153;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5153 (
            .in(out_5152),
            .outp(out_5153)
        );
        

        logic [WIDTH-1:0] out_5154;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5154 (
            .a(out_5150),
            .b(out_5153),
            .outp(out_5154)
        );        
        

        logic [WIDTH-1:0] out_5155;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5155 (
            .a(out_5144),
            .b(out_5154),
            .outp(out_5155)
        );        
        

        logic [WIDTH-1:0] out_5156;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.15)
        ) inst_5156 (
            .outp(out_5156)
        );
        

        logic [WIDTH-1:0] out_5157;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5157 (
            .a(out_14),
            .b(out_5156),
            .outp(out_5157)
        );        
        

        logic [WIDTH-1:0] out_5158;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5158 (
            .a(out_5153),
            .b(out_5157),
            .outp(out_5158)
        );        
        

        logic [WIDTH-1:0] out_5159;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5159 (
            .a(out_4929),
            .b(out_14),
            .outp(out_5159)
        );        
        

        logic [WIDTH-1:0] out_5160;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5160 (
            .a(out_5158),
            .b(out_5159),
            .outp(out_5160)
        );        
        

        logic [WIDTH-1:0] out_5161;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.72)
        ) inst_5161 (
            .outp(out_5161)
        );
        

        logic [WIDTH-1:0] out_5162;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5162 (
            .a(out_5161),
            .b(out_3),
            .outp(out_5162)
        );        
        

        logic [WIDTH-1:0] out_5163;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5163 (
            .a(out_5160),
            .b(out_5162),
            .outp(out_5163)
        );        
        

        logic [WIDTH-1:0] out_5164;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5164 (
            .in(out_4930),
            .outp(out_5164)
        );
        

        logic [WIDTH-1:0] out_5165;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.945)
        ) inst_5165 (
            .outp(out_5165)
        );
        

        logic [WIDTH-1:0] out_5166;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5166 (
            .a(out_5165),
            .b(out_3),
            .outp(out_5166)
        );        
        

        logic [WIDTH-1:0] out_5167;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5167 (
            .in(out_5166),
            .outp(out_5167)
        );
        

        logic [WIDTH-1:0] out_5168;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5168 (
            .a(out_5164),
            .b(out_5167),
            .outp(out_5168)
        );        
        

        logic [WIDTH-1:0] out_5169;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5169 (
            .in(out_5168),
            .outp(out_5169)
        );
        

        logic [WIDTH-1:0] out_5170;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5170 (
            .a(out_460),
            .b(out_5169),
            .outp(out_5170)
        );        
        

        logic [WIDTH-1:0] out_5171;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5171 (
            .a(out_5169),
            .b(out_9),
            .outp(out_5171)
        );        
        

        logic [WIDTH-1:0] out_5172;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5172 (
            .a(out_5170),
            .b(out_5171),
            .outp(out_5172)
        );        
        

        logic [WIDTH-1:0] out_5173;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.195)
        ) inst_5173 (
            .outp(out_5173)
        );
        

        logic [WIDTH-1:0] out_5174;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5174 (
            .a(out_5173),
            .b(out_3),
            .outp(out_5174)
        );        
        

        logic [WIDTH-1:0] out_5175;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5175 (
            .in(out_5174),
            .outp(out_5175)
        );
        

        logic [WIDTH-1:0] out_5176;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5176 (
            .a(out_5164),
            .b(out_5175),
            .outp(out_5176)
        );        
        

        logic [WIDTH-1:0] out_5177;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5177 (
            .in(out_5176),
            .outp(out_5177)
        );
        

        logic [WIDTH-1:0] out_5178;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5178 (
            .a(out_460),
            .b(out_5177),
            .outp(out_5178)
        );        
        

        logic [WIDTH-1:0] out_5179;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5179 (
            .a(out_5177),
            .b(out_9),
            .outp(out_5179)
        );        
        

        logic [WIDTH-1:0] out_5180;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5180 (
            .a(out_5178),
            .b(out_5179),
            .outp(out_5180)
        );        
        

        logic [WIDTH-1:0] out_5181;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5181 (
            .a(out_5172),
            .b(out_5180),
            .outp(out_5181)
        );        
        

        logic [WIDTH-1:0] out_5182;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5182 (
            .a(out_5163),
            .b(out_5181),
            .outp(out_5182)
        );        
        

        logic [WIDTH-1:0] out_5183;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5183 (
            .a(out_5155),
            .b(out_5182),
            .outp(out_5183)
        );        
        

        logic [WIDTH-1:0] out_5184;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.195)
        ) inst_5184 (
            .outp(out_5184)
        );
        

        logic [WIDTH-1:0] out_5185;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5185 (
            .a(out_5184),
            .b(out_152),
            .outp(out_5185)
        );        
        

        logic [WIDTH-1:0] out_5186;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.42975)
        ) inst_5186 (
            .outp(out_5186)
        );
        

        logic [WIDTH-1:0] out_5187;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5187 (
            .a(out_5186),
            .b(out_127),
            .outp(out_5187)
        );        
        

        logic [WIDTH-1:0] out_5188;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5188 (
            .a(out_5187),
            .b(out_1011),
            .outp(out_5188)
        );        
        

        logic [WIDTH-1:0] out_5189;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5189 (
            .a(out_5185),
            .b(out_5188),
            .outp(out_5189)
        );        
        

        logic [WIDTH-1:0] out_5190;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.67975)
        ) inst_5190 (
            .outp(out_5190)
        );
        

        logic [WIDTH-1:0] out_5191;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5191 (
            .a(out_5190),
            .b(out_127),
            .outp(out_5191)
        );        
        

        logic [WIDTH-1:0] out_5192;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5192 (
            .a(out_1017),
            .b(out_5191),
            .outp(out_5192)
        );        
        

        logic [WIDTH-1:0] out_5193;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5193 (
            .a(out_5189),
            .b(out_5192),
            .outp(out_5193)
        );        
        

        logic [WIDTH-1:0] out_5194;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5194 (
            .a(out_5183),
            .b(out_5193),
            .outp(out_5194)
        );        
        

        logic [WIDTH-1:0] out_5195;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5195 (
            .a(out_5191),
            .b(out_1017),
            .outp(out_5195)
        );        
        

        logic [WIDTH-1:0] out_5196;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5196 (
            .a(out_1011),
            .b(out_5187),
            .outp(out_5196)
        );        
        

        logic [WIDTH-1:0] out_5197;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5197 (
            .a(out_5195),
            .b(out_5196),
            .outp(out_5197)
        );        
        

        logic [WIDTH-1:0] out_5198;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5198 (
            .a(out_152),
            .b(out_5184),
            .outp(out_5198)
        );        
        

        logic [WIDTH-1:0] out_5199;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5199 (
            .a(out_5197),
            .b(out_5198),
            .outp(out_5199)
        );        
        

        logic [WIDTH-1:0] out_5200;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5200 (
            .a(out_5194),
            .b(out_5199),
            .outp(out_5200)
        );        
        

        logic [WIDTH-1:0] out_5201;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.25)
        ) inst_5201 (
            .outp(out_5201)
        );
        

        logic [WIDTH-1:0] out_5202;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5202 (
            .a(out_137),
            .b(out_5201),
            .outp(out_5202)
        );        
        

        logic [WIDTH-1:0] out_5203;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5203 (
            .a(out_5195),
            .b(out_5202),
            .outp(out_5203)
        );        
        

        logic [WIDTH-1:0] out_5204;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.48475)
        ) inst_5204 (
            .outp(out_5204)
        );
        

        logic [WIDTH-1:0] out_5205;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5205 (
            .a(out_5204),
            .b(out_127),
            .outp(out_5205)
        );        
        

        logic [WIDTH-1:0] out_5206;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5206 (
            .a(out_1011),
            .b(out_5205),
            .outp(out_5206)
        );        
        

        logic [WIDTH-1:0] out_5207;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5207 (
            .a(out_5203),
            .b(out_5206),
            .outp(out_5207)
        );        
        

        logic [WIDTH-1:0] out_5208;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5208 (
            .a(out_5200),
            .b(out_5207),
            .outp(out_5208)
        );        
        

        logic [WIDTH-1:0] out_5209;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5209 (
            .a(out_5205),
            .b(out_1011),
            .outp(out_5209)
        );        
        

        logic [WIDTH-1:0] out_5210;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5210 (
            .a(out_5192),
            .b(out_5209),
            .outp(out_5210)
        );        
        

        logic [WIDTH-1:0] out_5211;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5211 (
            .a(out_5201),
            .b(out_137),
            .outp(out_5211)
        );        
        

        logic [WIDTH-1:0] out_5212;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5212 (
            .a(out_5210),
            .b(out_5211),
            .outp(out_5212)
        );        
        

        logic [WIDTH-1:0] out_5213;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5213 (
            .a(out_5208),
            .b(out_5212),
            .outp(out_5213)
        );        
        

        logic [WIDTH-1:0] out_5214;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5214 (
            .a(out_4447),
            .b(out_5188),
            .outp(out_5214)
        );        
        

        logic [WIDTH-1:0] out_5215;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.73475)
        ) inst_5215 (
            .outp(out_5215)
        );
        

        logic [WIDTH-1:0] out_5216;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5216 (
            .a(out_5215),
            .b(out_127),
            .outp(out_5216)
        );        
        

        logic [WIDTH-1:0] out_5217;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5217 (
            .a(out_1017),
            .b(out_5216),
            .outp(out_5217)
        );        
        

        logic [WIDTH-1:0] out_5218;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5218 (
            .a(out_5214),
            .b(out_5217),
            .outp(out_5218)
        );        
        

        logic [WIDTH-1:0] out_5219;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5219 (
            .a(out_5213),
            .b(out_5218),
            .outp(out_5219)
        );        
        

        logic [WIDTH-1:0] out_5220;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5220 (
            .a(out_4460),
            .b(out_5196),
            .outp(out_5220)
        );        
        

        logic [WIDTH-1:0] out_5221;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5221 (
            .a(out_5216),
            .b(out_1017),
            .outp(out_5221)
        );        
        

        logic [WIDTH-1:0] out_5222;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5222 (
            .a(out_5220),
            .b(out_5221),
            .outp(out_5222)
        );        
        

        logic [WIDTH-1:0] out_5223;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5223 (
            .a(out_5219),
            .b(out_5222),
            .outp(out_5223)
        );        
        

        logic [WIDTH-1:0] out_5224;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5224 (
            .a(out_4464),
            .b(out_5206),
            .outp(out_5224)
        );        
        

        logic [WIDTH-1:0] out_5225;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5225 (
            .a(out_5224),
            .b(out_5221),
            .outp(out_5225)
        );        
        

        logic [WIDTH-1:0] out_5226;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5226 (
            .a(out_5223),
            .b(out_5225),
            .outp(out_5226)
        );        
        

        logic [WIDTH-1:0] out_5227;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5227 (
            .a(out_4473),
            .b(out_5209),
            .outp(out_5227)
        );        
        

        logic [WIDTH-1:0] out_5228;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5228 (
            .a(out_5227),
            .b(out_5217),
            .outp(out_5228)
        );        
        

        logic [WIDTH-1:0] out_5229;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5229 (
            .a(out_5226),
            .b(out_5228),
            .outp(out_5229)
        );        
        

        logic [WIDTH-1:0] out_5230;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.35975)
        ) inst_5230 (
            .outp(out_5230)
        );
        

        logic [WIDTH-1:0] out_5231;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5231 (
            .a(out_5230),
            .b(out_1011),
            .outp(out_5231)
        );        
        

        logic [WIDTH-1:0] out_5232;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5232 (
            .a(out_5231),
            .b(out_127),
            .outp(out_5232)
        );        
        

        logic [WIDTH-1:0] out_5233;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5233 (
            .in(out_5232),
            .outp(out_5233)
        );
        

        logic [WIDTH-1:0] out_5234;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5234 (
            .a(out_4447),
            .b(out_5233),
            .outp(out_5234)
        );        
        

        logic [WIDTH-1:0] out_5235;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.05475)
        ) inst_5235 (
            .outp(out_5235)
        );
        

        logic [WIDTH-1:0] out_5236;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5236 (
            .a(out_5235),
            .b(out_1017),
            .outp(out_5236)
        );        
        

        logic [WIDTH-1:0] out_5237;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5237 (
            .a(out_5236),
            .b(out_127),
            .outp(out_5237)
        );        
        

        logic [WIDTH-1:0] out_5238;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5238 (
            .a(out_5234),
            .b(out_5237),
            .outp(out_5238)
        );        
        

        logic [WIDTH-1:0] out_5239;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5239 (
            .a(out_5229),
            .b(out_5238),
            .outp(out_5239)
        );        
        

        logic [WIDTH-1:0] out_5240;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5240 (
            .a(out_4460),
            .b(out_5232),
            .outp(out_5240)
        );        
        

        logic [WIDTH-1:0] out_5241;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5241 (
            .in(out_5237),
            .outp(out_5241)
        );
        

        logic [WIDTH-1:0] out_5242;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5242 (
            .a(out_5240),
            .b(out_5241),
            .outp(out_5242)
        );        
        

        logic [WIDTH-1:0] out_5243;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5243 (
            .a(out_5239),
            .b(out_5242),
            .outp(out_5243)
        );        
        

        logic [WIDTH-1:0] out_5244;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5244 (
            .a(out_4464),
            .b(out_5241),
            .outp(out_5244)
        );        
        

        logic [WIDTH-1:0] out_5245;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.30475)
        ) inst_5245 (
            .outp(out_5245)
        );
        

        logic [WIDTH-1:0] out_5246;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5246 (
            .a(out_5245),
            .b(out_1011),
            .outp(out_5246)
        );        
        

        logic [WIDTH-1:0] out_5247;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5247 (
            .a(out_5246),
            .b(out_127),
            .outp(out_5247)
        );        
        

        logic [WIDTH-1:0] out_5248;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5248 (
            .a(out_5244),
            .b(out_5247),
            .outp(out_5248)
        );        
        

        logic [WIDTH-1:0] out_5249;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5249 (
            .a(out_5243),
            .b(out_5248),
            .outp(out_5249)
        );        
        

        logic [WIDTH-1:0] out_5250;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5250 (
            .a(out_4473),
            .b(out_5237),
            .outp(out_5250)
        );        
        

        logic [WIDTH-1:0] out_5251;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5251 (
            .in(out_5247),
            .outp(out_5251)
        );
        

        logic [WIDTH-1:0] out_5252;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5252 (
            .a(out_5250),
            .b(out_5251),
            .outp(out_5252)
        );        
        

        logic [WIDTH-1:0] out_5253;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5253 (
            .a(out_5249),
            .b(out_5252),
            .outp(out_5253)
        );        
        

        logic [WIDTH-1:0] out_5254;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.725)
        ) inst_5254 (
            .outp(out_5254)
        );
        

        logic [WIDTH-1:0] out_5255;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5255 (
            .a(out_5254),
            .b(out_3),
            .outp(out_5255)
        );        
        

        logic [WIDTH-1:0] out_5256;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5256 (
            .in(out_5255),
            .outp(out_5256)
        );
        

        logic [WIDTH-1:0] out_5257;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5257 (
            .a(out_3384),
            .b(out_5256),
            .outp(out_5257)
        );        
        

        logic [WIDTH-1:0] out_5258;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0749998)
        ) inst_5258 (
            .outp(out_5258)
        );
        

        logic [WIDTH-1:0] out_5259;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5259 (
            .a(out_5258),
            .b(out_14),
            .outp(out_5259)
        );        
        

        logic [WIDTH-1:0] out_5260;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5260 (
            .in(out_5259),
            .outp(out_5260)
        );
        

        logic [WIDTH-1:0] out_5261;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5261 (
            .a(out_5257),
            .b(out_5260),
            .outp(out_5261)
        );        
        

        logic [WIDTH-1:0] out_5262;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.625)
        ) inst_5262 (
            .outp(out_5262)
        );
        

        logic [WIDTH-1:0] out_5263;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5263 (
            .a(out_5262),
            .b(out_3),
            .outp(out_5263)
        );        
        

        logic [WIDTH-1:0] out_5264;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5264 (
            .a(out_5261),
            .b(out_5263),
            .outp(out_5264)
        );        
        

        logic [WIDTH-1:0] out_5265;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5265 (
            .a(out_5253),
            .b(out_5264),
            .outp(out_5265)
        );        
        

        logic [WIDTH-1:0] out_5266;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.45)
        ) inst_5266 (
            .outp(out_5266)
        );
        

        logic [WIDTH-1:0] out_5267;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5267 (
            .a(out_5266),
            .b(out_3),
            .outp(out_5267)
        );        
        

        logic [WIDTH-1:0] out_5268;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5268 (
            .in(out_5267),
            .outp(out_5268)
        );
        

        logic [WIDTH-1:0] out_5269;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5269 (
            .a(out_3147),
            .b(out_5268),
            .outp(out_5269)
        );        
        

        logic [WIDTH-1:0] out_5270;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5270 (
            .in(out_5269),
            .outp(out_5270)
        );
        

        logic [WIDTH-1:0] out_5271;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5271 (
            .a(out_9),
            .b(out_5270),
            .outp(out_5271)
        );        
        

        logic [WIDTH-1:0] out_5272;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5272 (
            .a(out_5270),
            .b(out_21),
            .outp(out_5272)
        );        
        

        logic [WIDTH-1:0] out_5273;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5273 (
            .a(out_5271),
            .b(out_5272),
            .outp(out_5273)
        );        
        

        logic [WIDTH-1:0] out_5274;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5274 (
            .a(out_5265),
            .b(out_5273),
            .outp(out_5274)
        );        
        

        logic [WIDTH-1:0] out_5275;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.825)
        ) inst_5275 (
            .outp(out_5275)
        );
        

        logic [WIDTH-1:0] out_5276;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5276 (
            .a(out_5275),
            .b(out_3),
            .outp(out_5276)
        );        
        

        logic [WIDTH-1:0] out_5277;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5277 (
            .a(out_3464),
            .b(out_5276),
            .outp(out_5277)
        );        
        

        logic [WIDTH-1:0] out_5278;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5278 (
            .in(out_685),
            .outp(out_5278)
        );
        

        logic [WIDTH-1:0] out_5279;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5279 (
            .a(out_5277),
            .b(out_5278),
            .outp(out_5279)
        );        
        

        logic [WIDTH-1:0] out_5280;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5280 (
            .a(out_5274),
            .b(out_5279),
            .outp(out_5280)
        );        
        

        logic [WIDTH-1:0] out_5281;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5281 (
            .a(out_3384),
            .b(out_3386),
            .outp(out_5281)
        );        
        

        logic [WIDTH-1:0] out_5282;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.275)
        ) inst_5282 (
            .outp(out_5282)
        );
        

        logic [WIDTH-1:0] out_5283;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5283 (
            .a(out_5282),
            .b(out_3),
            .outp(out_5283)
        );        
        

        logic [WIDTH-1:0] out_5284;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5284 (
            .a(out_5281),
            .b(out_5283),
            .outp(out_5284)
        );        
        

        logic [WIDTH-1:0] out_5285;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.375)
        ) inst_5285 (
            .outp(out_5285)
        );
        

        logic [WIDTH-1:0] out_5286;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5286 (
            .a(out_5285),
            .b(out_3),
            .outp(out_5286)
        );        
        

        logic [WIDTH-1:0] out_5287;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5287 (
            .in(out_5286),
            .outp(out_5287)
        );
        

        logic [WIDTH-1:0] out_5288;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5288 (
            .a(out_5284),
            .b(out_5287),
            .outp(out_5288)
        );        
        

        logic [WIDTH-1:0] out_5289;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5289 (
            .a(out_5280),
            .b(out_5288),
            .outp(out_5289)
        );        
        

        logic [WIDTH-1:0] out_5290;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5290 (
            .a(out_3366),
            .b(out_5276),
            .outp(out_5290)
        );        
        

        logic [WIDTH-1:0] out_5291;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5291 (
            .a(out_5290),
            .b(out_5287),
            .outp(out_5291)
        );        
        

        logic [WIDTH-1:0] out_5292;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.1)
        ) inst_5292 (
            .outp(out_5292)
        );
        

        logic [WIDTH-1:0] out_5293;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5293 (
            .a(out_5292),
            .b(out_3),
            .outp(out_5293)
        );        
        

        logic [WIDTH-1:0] out_5294;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5294 (
            .in(out_5293),
            .outp(out_5294)
        );
        

        logic [WIDTH-1:0] out_5295;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5295 (
            .a(out_3147),
            .b(out_5294),
            .outp(out_5295)
        );        
        

        logic [WIDTH-1:0] out_5296;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5296 (
            .in(out_5295),
            .outp(out_5296)
        );
        

        logic [WIDTH-1:0] out_5297;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5297 (
            .a(out_9),
            .b(out_5296),
            .outp(out_5297)
        );        
        

        logic [WIDTH-1:0] out_5298;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5298 (
            .a(out_5291),
            .b(out_5297),
            .outp(out_5298)
        );        
        

        logic [WIDTH-1:0] out_5299;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5299 (
            .a(out_5296),
            .b(out_21),
            .outp(out_5299)
        );        
        

        logic [WIDTH-1:0] out_5300;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5300 (
            .a(out_5298),
            .b(out_5299),
            .outp(out_5300)
        );        
        

        logic [WIDTH-1:0] out_5301;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5301 (
            .a(out_5289),
            .b(out_5300),
            .outp(out_5301)
        );        
        

        logic [WIDTH-1:0] out_5302;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.275)
        ) inst_5302 (
            .outp(out_5302)
        );
        

        logic [WIDTH-1:0] out_5303;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5303 (
            .a(out_5302),
            .b(out_3),
            .outp(out_5303)
        );        
        

        logic [WIDTH-1:0] out_5304;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5304 (
            .in(out_5303),
            .outp(out_5304)
        );
        

        logic [WIDTH-1:0] out_5305;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5305 (
            .a(out_3374),
            .b(out_5304),
            .outp(out_5305)
        );        
        

        logic [WIDTH-1:0] out_5306;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.175)
        ) inst_5306 (
            .outp(out_5306)
        );
        

        logic [WIDTH-1:0] out_5307;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5307 (
            .a(out_5306),
            .b(out_3),
            .outp(out_5307)
        );        
        

        logic [WIDTH-1:0] out_5308;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5308 (
            .a(out_5305),
            .b(out_5307),
            .outp(out_5308)
        );        
        

        logic [WIDTH-1:0] out_5309;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5309 (
            .a(out_5301),
            .b(out_5308),
            .outp(out_5309)
        );        
        

        logic [WIDTH-1:0] out_5310;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.75)
        ) inst_5310 (
            .outp(out_5310)
        );
        

        logic [WIDTH-1:0] out_5311;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5311 (
            .a(out_5310),
            .b(out_14),
            .outp(out_5311)
        );        
        

        logic [WIDTH-1:0] out_5312;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5312 (
            .a(out_3384),
            .b(out_5311),
            .outp(out_5312)
        );        
        

        logic [WIDTH-1:0] out_5313;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.45)
        ) inst_5313 (
            .outp(out_5313)
        );
        

        logic [WIDTH-1:0] out_5314;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5314 (
            .a(out_5313),
            .b(out_3),
            .outp(out_5314)
        );        
        

        logic [WIDTH-1:0] out_5315;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5315 (
            .in(out_5314),
            .outp(out_5315)
        );
        

        logic [WIDTH-1:0] out_5316;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5316 (
            .a(out_5312),
            .b(out_5315),
            .outp(out_5316)
        );        
        

        logic [WIDTH-1:0] out_5317;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.275)
        ) inst_5317 (
            .outp(out_5317)
        );
        

        logic [WIDTH-1:0] out_5318;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5318 (
            .a(out_5317),
            .b(out_3),
            .outp(out_5318)
        );        
        

        logic [WIDTH-1:0] out_5319;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5319 (
            .a(out_5316),
            .b(out_5318),
            .outp(out_5319)
        );        
        

        logic [WIDTH-1:0] out_5320;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5320 (
            .a(out_5309),
            .b(out_5319),
            .outp(out_5320)
        );        
        

        logic [WIDTH-1:0] out_5321;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5321 (
            .a(out_3124),
            .b(out_5315),
            .outp(out_5321)
        );        
        

        logic [WIDTH-1:0] out_5322;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5322 (
            .a(out_5321),
            .b(out_5318),
            .outp(out_5322)
        );        
        

        logic [WIDTH-1:0] out_5323;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4)
        ) inst_5323 (
            .outp(out_5323)
        );
        

        logic [WIDTH-1:0] out_5324;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5324 (
            .a(out_14),
            .b(out_5323),
            .outp(out_5324)
        );        
        

        logic [WIDTH-1:0] out_5325;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5325 (
            .a(out_5322),
            .b(out_5324),
            .outp(out_5325)
        );        
        

        logic [WIDTH-1:0] out_5326;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5326 (
            .a(out_5320),
            .b(out_5325),
            .outp(out_5326)
        );        
        

        logic [WIDTH-1:0] out_5327;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5327 (
            .a(out_3374),
            .b(out_5314),
            .outp(out_5327)
        );        
        

        logic [WIDTH-1:0] out_5328;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.175)
        ) inst_5328 (
            .outp(out_5328)
        );
        

        logic [WIDTH-1:0] out_5329;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5329 (
            .a(out_5328),
            .b(out_3),
            .outp(out_5329)
        );        
        

        logic [WIDTH-1:0] out_5330;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5330 (
            .in(out_5329),
            .outp(out_5330)
        );
        

        logic [WIDTH-1:0] out_5331;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5331 (
            .a(out_5327),
            .b(out_5330),
            .outp(out_5331)
        );        
        

        logic [WIDTH-1:0] out_5332;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5332 (
            .in(out_5315),
            .outp(out_5332)
        );
        

        logic [WIDTH-1:0] out_5333;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5333 (
            .a(out_3147),
            .b(out_5332),
            .outp(out_5333)
        );        
        

        logic [WIDTH-1:0] out_5334;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5334 (
            .in(out_5333),
            .outp(out_5334)
        );
        

        logic [WIDTH-1:0] out_5335;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5335 (
            .a(out_9),
            .b(out_5334),
            .outp(out_5335)
        );        
        

        logic [WIDTH-1:0] out_5336;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5336 (
            .a(out_5331),
            .b(out_5335),
            .outp(out_5336)
        );        
        

        logic [WIDTH-1:0] out_5337;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5337 (
            .a(out_5334),
            .b(out_21),
            .outp(out_5337)
        );        
        

        logic [WIDTH-1:0] out_5338;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5338 (
            .a(out_5336),
            .b(out_5337),
            .outp(out_5338)
        );        
        

        logic [WIDTH-1:0] out_5339;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5339 (
            .a(out_5326),
            .b(out_5338),
            .outp(out_5339)
        );        
        

        logic [WIDTH-1:0] out_5340;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5340 (
            .a(out_3124),
            .b(out_3044),
            .outp(out_5340)
        );        
        

        logic [WIDTH-1:0] out_5341;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5341 (
            .a(out_5340),
            .b(out_3275),
            .outp(out_5341)
        );        
        

        logic [WIDTH-1:0] out_5342;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5342 (
            .in(out_3071),
            .outp(out_5342)
        );
        

        logic [WIDTH-1:0] out_5343;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5343 (
            .a(out_5341),
            .b(out_5342),
            .outp(out_5343)
        );        
        

        logic [WIDTH-1:0] out_5344;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5344 (
            .a(out_5339),
            .b(out_5343),
            .outp(out_5344)
        );        
        

        logic [WIDTH-1:0] out_5345;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.25)
        ) inst_5345 (
            .outp(out_5345)
        );
        

        logic [WIDTH-1:0] out_5346;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5346 (
            .a(out_5345),
            .b(out_3),
            .outp(out_5346)
        );        
        

        logic [WIDTH-1:0] out_5347;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5347 (
            .a(out_3464),
            .b(out_5346),
            .outp(out_5347)
        );        
        

        logic [WIDTH-1:0] out_5348;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.35)
        ) inst_5348 (
            .outp(out_5348)
        );
        

        logic [WIDTH-1:0] out_5349;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5349 (
            .a(out_5348),
            .b(out_3),
            .outp(out_5349)
        );        
        

        logic [WIDTH-1:0] out_5350;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5350 (
            .in(out_5349),
            .outp(out_5350)
        );
        

        logic [WIDTH-1:0] out_5351;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5351 (
            .a(out_5347),
            .b(out_5350),
            .outp(out_5351)
        );        
        

        logic [WIDTH-1:0] out_5352;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5352 (
            .a(out_5344),
            .b(out_5351),
            .outp(out_5352)
        );        
        

        logic [WIDTH-1:0] out_5353;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.025)
        ) inst_5353 (
            .outp(out_5353)
        );
        

        logic [WIDTH-1:0] out_5354;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5354 (
            .a(out_5353),
            .b(out_3),
            .outp(out_5354)
        );        
        

        logic [WIDTH-1:0] out_5355;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5355 (
            .a(out_3366),
            .b(out_5354),
            .outp(out_5355)
        );        
        

        logic [WIDTH-1:0] out_5356;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.125)
        ) inst_5356 (
            .outp(out_5356)
        );
        

        logic [WIDTH-1:0] out_5357;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5357 (
            .a(out_5356),
            .b(out_3),
            .outp(out_5357)
        );        
        

        logic [WIDTH-1:0] out_5358;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5358 (
            .in(out_5357),
            .outp(out_5358)
        );
        

        logic [WIDTH-1:0] out_5359;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5359 (
            .a(out_5355),
            .b(out_5358),
            .outp(out_5359)
        );        
        

        logic [WIDTH-1:0] out_5360;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5360 (
            .a(out_5352),
            .b(out_5359),
            .outp(out_5360)
        );        
        

        logic [WIDTH-1:0] out_5361;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.475)
        ) inst_5361 (
            .outp(out_5361)
        );
        

        logic [WIDTH-1:0] out_5362;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5362 (
            .a(out_5361),
            .b(out_3),
            .outp(out_5362)
        );        
        

        logic [WIDTH-1:0] out_5363;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5363 (
            .a(out_3374),
            .b(out_5362),
            .outp(out_5363)
        );        
        

        logic [WIDTH-1:0] out_5364;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.575)
        ) inst_5364 (
            .outp(out_5364)
        );
        

        logic [WIDTH-1:0] out_5365;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5365 (
            .a(out_5364),
            .b(out_3),
            .outp(out_5365)
        );        
        

        logic [WIDTH-1:0] out_5366;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5366 (
            .in(out_5365),
            .outp(out_5366)
        );
        

        logic [WIDTH-1:0] out_5367;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5367 (
            .a(out_5363),
            .b(out_5366),
            .outp(out_5367)
        );        
        

        logic [WIDTH-1:0] out_5368;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5368 (
            .a(out_5360),
            .b(out_5367),
            .outp(out_5368)
        );        
        

        logic [WIDTH-1:0] out_5369;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5369 (
            .a(out_5281),
            .b(out_5354),
            .outp(out_5369)
        );        
        

        logic [WIDTH-1:0] out_5370;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5370 (
            .a(out_5369),
            .b(out_5366),
            .outp(out_5370)
        );        
        

        logic [WIDTH-1:0] out_5371;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5371 (
            .a(out_3096),
            .b(out_3),
            .outp(out_5371)
        );        
        

        logic [WIDTH-1:0] out_5372;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5372 (
            .in(out_5371),
            .outp(out_5372)
        );
        

        logic [WIDTH-1:0] out_5373;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5373 (
            .a(out_3147),
            .b(out_5372),
            .outp(out_5373)
        );        
        

        logic [WIDTH-1:0] out_5374;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5374 (
            .in(out_5373),
            .outp(out_5374)
        );
        

        logic [WIDTH-1:0] out_5375;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5375 (
            .a(out_9),
            .b(out_5374),
            .outp(out_5375)
        );        
        

        logic [WIDTH-1:0] out_5376;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5376 (
            .a(out_5370),
            .b(out_5375),
            .outp(out_5376)
        );        
        

        logic [WIDTH-1:0] out_5377;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5377 (
            .a(out_5374),
            .b(out_21),
            .outp(out_5377)
        );        
        

        logic [WIDTH-1:0] out_5378;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5378 (
            .a(out_5376),
            .b(out_5377),
            .outp(out_5378)
        );        
        

        logic [WIDTH-1:0] out_5379;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5379 (
            .a(out_5368),
            .b(out_5378),
            .outp(out_5379)
        );        
        

        logic [WIDTH-1:0] out_5380;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.825)
        ) inst_5380 (
            .outp(out_5380)
        );
        

        logic [WIDTH-1:0] out_5381;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5381 (
            .a(out_5380),
            .b(out_3),
            .outp(out_5381)
        );        
        

        logic [WIDTH-1:0] out_5382;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5382 (
            .a(out_3100),
            .b(out_5381),
            .outp(out_5382)
        );        
        

        logic [WIDTH-1:0] out_5383;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.925)
        ) inst_5383 (
            .outp(out_5383)
        );
        

        logic [WIDTH-1:0] out_5384;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5384 (
            .a(out_5383),
            .b(out_3),
            .outp(out_5384)
        );        
        

        logic [WIDTH-1:0] out_5385;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5385 (
            .in(out_5384),
            .outp(out_5385)
        );
        

        logic [WIDTH-1:0] out_5386;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5386 (
            .a(out_5382),
            .b(out_5385),
            .outp(out_5386)
        );        
        

        logic [WIDTH-1:0] out_5387;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5387 (
            .a(out_5379),
            .b(out_5386),
            .outp(out_5387)
        );        
        

        logic [WIDTH-1:0] out_5388;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5388 (
            .a(out_4532),
            .b(out_3),
            .outp(out_5388)
        );        
        

        logic [WIDTH-1:0] out_5389;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5389 (
            .a(out_3112),
            .b(out_5388),
            .outp(out_5389)
        );        
        

        logic [WIDTH-1:0] out_5390;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.075)
        ) inst_5390 (
            .outp(out_5390)
        );
        

        logic [WIDTH-1:0] out_5391;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5391 (
            .a(out_5390),
            .b(out_3),
            .outp(out_5391)
        );        
        

        logic [WIDTH-1:0] out_5392;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5392 (
            .in(out_5391),
            .outp(out_5392)
        );
        

        logic [WIDTH-1:0] out_5393;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5393 (
            .a(out_5389),
            .b(out_5392),
            .outp(out_5393)
        );        
        

        logic [WIDTH-1:0] out_5394;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5394 (
            .a(out_5387),
            .b(out_5393),
            .outp(out_5394)
        );        
        

        logic [WIDTH-1:0] out_5395;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5395 (
            .a(out_3412),
            .b(out_5388),
            .outp(out_5395)
        );        
        

        logic [WIDTH-1:0] out_5396;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5396 (
            .a(out_5395),
            .b(out_5392),
            .outp(out_5396)
        );        
        

        logic [WIDTH-1:0] out_5397;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5397 (
            .in(out_5388),
            .outp(out_5397)
        );
        

        logic [WIDTH-1:0] out_5398;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5398 (
            .a(out_3126),
            .b(out_5397),
            .outp(out_5398)
        );        
        

        logic [WIDTH-1:0] out_5399;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5399 (
            .in(out_5398),
            .outp(out_5399)
        );
        

        logic [WIDTH-1:0] out_5400;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5400 (
            .a(out_336),
            .b(out_5399),
            .outp(out_5400)
        );        
        

        logic [WIDTH-1:0] out_5401;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5401 (
            .a(out_5396),
            .b(out_5400),
            .outp(out_5401)
        );        
        

        logic [WIDTH-1:0] out_5402;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5402 (
            .a(out_5399),
            .b(out_343),
            .outp(out_5402)
        );        
        

        logic [WIDTH-1:0] out_5403;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5403 (
            .a(out_5401),
            .b(out_5402),
            .outp(out_5403)
        );        
        

        logic [WIDTH-1:0] out_5404;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5404 (
            .a(out_5394),
            .b(out_5403),
            .outp(out_5404)
        );        
        

        logic [WIDTH-1:0] out_5405;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.875)
        ) inst_5405 (
            .outp(out_5405)
        );
        

        logic [WIDTH-1:0] out_5406;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5406 (
            .a(out_5405),
            .b(out_3),
            .outp(out_5406)
        );        
        

        logic [WIDTH-1:0] out_5407;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5407 (
            .a(out_3564),
            .b(out_5406),
            .outp(out_5407)
        );        
        

        logic [WIDTH-1:0] out_5408;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.975)
        ) inst_5408 (
            .outp(out_5408)
        );
        

        logic [WIDTH-1:0] out_5409;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5409 (
            .a(out_5408),
            .b(out_3),
            .outp(out_5409)
        );        
        

        logic [WIDTH-1:0] out_5410;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5410 (
            .in(out_5409),
            .outp(out_5410)
        );
        

        logic [WIDTH-1:0] out_5411;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5411 (
            .a(out_5407),
            .b(out_5410),
            .outp(out_5411)
        );        
        

        logic [WIDTH-1:0] out_5412;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5412 (
            .a(out_5404),
            .b(out_5411),
            .outp(out_5412)
        );        
        

        logic [WIDTH-1:0] out_5413;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.325)
        ) inst_5413 (
            .outp(out_5413)
        );
        

        logic [WIDTH-1:0] out_5414;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5414 (
            .a(out_5413),
            .b(out_3),
            .outp(out_5414)
        );        
        

        logic [WIDTH-1:0] out_5415;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5415 (
            .a(out_3464),
            .b(out_5414),
            .outp(out_5415)
        );        
        

        logic [WIDTH-1:0] out_5416;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.425)
        ) inst_5416 (
            .outp(out_5416)
        );
        

        logic [WIDTH-1:0] out_5417;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5417 (
            .a(out_5416),
            .b(out_3),
            .outp(out_5417)
        );        
        

        logic [WIDTH-1:0] out_5418;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5418 (
            .in(out_5417),
            .outp(out_5418)
        );
        

        logic [WIDTH-1:0] out_5419;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5419 (
            .a(out_5415),
            .b(out_5418),
            .outp(out_5419)
        );        
        

        logic [WIDTH-1:0] out_5420;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5420 (
            .a(out_5412),
            .b(out_5419),
            .outp(out_5420)
        );        
        

        logic [WIDTH-1:0] out_5421;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5421 (
            .a(out_3384),
            .b(out_3582),
            .outp(out_5421)
        );        
        

        logic [WIDTH-1:0] out_5422;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5422 (
            .a(out_5421),
            .b(out_5406),
            .outp(out_5422)
        );        
        

        logic [WIDTH-1:0] out_5423;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5423 (
            .a(out_5422),
            .b(out_5418),
            .outp(out_5423)
        );        
        

        logic [WIDTH-1:0] out_5424;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5424 (
            .a(out_5156),
            .b(out_3),
            .outp(out_5424)
        );        
        

        logic [WIDTH-1:0] out_5425;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5425 (
            .in(out_5424),
            .outp(out_5425)
        );
        

        logic [WIDTH-1:0] out_5426;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5426 (
            .a(out_3147),
            .b(out_5425),
            .outp(out_5426)
        );        
        

        logic [WIDTH-1:0] out_5427;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5427 (
            .in(out_5426),
            .outp(out_5427)
        );
        

        logic [WIDTH-1:0] out_5428;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5428 (
            .a(out_9),
            .b(out_5427),
            .outp(out_5428)
        );        
        

        logic [WIDTH-1:0] out_5429;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5429 (
            .a(out_5423),
            .b(out_5428),
            .outp(out_5429)
        );        
        

        logic [WIDTH-1:0] out_5430;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5430 (
            .a(out_5427),
            .b(out_21),
            .outp(out_5430)
        );        
        

        logic [WIDTH-1:0] out_5431;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5431 (
            .a(out_5429),
            .b(out_5430),
            .outp(out_5431)
        );        
        

        logic [WIDTH-1:0] out_5432;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5432 (
            .a(out_5420),
            .b(out_5431),
            .outp(out_5432)
        );        
        

        logic [WIDTH-1:0] out_5433;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.8)
        ) inst_5433 (
            .outp(out_5433)
        );
        

        logic [WIDTH-1:0] out_5434;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5434 (
            .a(out_5433),
            .b(out_3),
            .outp(out_5434)
        );        
        

        logic [WIDTH-1:0] out_5435;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5435 (
            .in(out_5434),
            .outp(out_5435)
        );
        

        logic [WIDTH-1:0] out_5436;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5436 (
            .a(out_3147),
            .b(out_5435),
            .outp(out_5436)
        );        
        

        logic [WIDTH-1:0] out_5437;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5437 (
            .in(out_5436),
            .outp(out_5437)
        );
        

        logic [WIDTH-1:0] out_5438;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5438 (
            .a(out_9),
            .b(out_5437),
            .outp(out_5438)
        );        
        

        logic [WIDTH-1:0] out_5439;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5439 (
            .a(out_5437),
            .b(out_21),
            .outp(out_5439)
        );        
        

        logic [WIDTH-1:0] out_5440;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5440 (
            .a(out_5438),
            .b(out_5439),
            .outp(out_5440)
        );        
        

        logic [WIDTH-1:0] out_5441;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5441 (
            .a(out_5432),
            .b(out_5440),
            .outp(out_5441)
        );        
        

        logic [WIDTH-1:0] out_5442;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5442 (
            .a(out_4551),
            .b(out_4559),
            .outp(out_5442)
        );        
        

        logic [WIDTH-1:0] out_5443;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.958)
        ) inst_5443 (
            .outp(out_5443)
        );
        

        logic [WIDTH-1:0] out_5444;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5444 (
            .a(out_3),
            .b(out_5443),
            .outp(out_5444)
        );        
        

        logic [WIDTH-1:0] out_5445;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5445 (
            .a(out_5442),
            .b(out_5444),
            .outp(out_5445)
        );        
        

        logic [WIDTH-1:0] out_5446;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.858)
        ) inst_5446 (
            .outp(out_5446)
        );
        

        logic [WIDTH-1:0] out_5447;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5447 (
            .a(out_5446),
            .b(out_3),
            .outp(out_5447)
        );        
        

        logic [WIDTH-1:0] out_5448;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5448 (
            .a(out_5445),
            .b(out_5447),
            .outp(out_5448)
        );        
        

        logic [WIDTH-1:0] out_5449;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5449 (
            .a(out_5441),
            .b(out_5448),
            .outp(out_5449)
        );        
        

        logic [WIDTH-1:0] out_5450;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.133)
        ) inst_5450 (
            .outp(out_5450)
        );
        

        logic [WIDTH-1:0] out_5451;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5451 (
            .a(out_3),
            .b(out_5450),
            .outp(out_5451)
        );        
        

        logic [WIDTH-1:0] out_5452;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5452 (
            .in(out_5451),
            .outp(out_5452)
        );
        

        logic [WIDTH-1:0] out_5453;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5453 (
            .a(out_5452),
            .b(out_4534),
            .outp(out_5453)
        );        
        

        logic [WIDTH-1:0] out_5454;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5454 (
            .in(out_5453),
            .outp(out_5454)
        );
        

        logic [WIDTH-1:0] out_5455;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5455 (
            .a(out_9),
            .b(out_5454),
            .outp(out_5455)
        );        
        

        logic [WIDTH-1:0] out_5456;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5456 (
            .a(out_4573),
            .b(out_5455),
            .outp(out_5456)
        );        
        

        logic [WIDTH-1:0] out_5457;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5457 (
            .a(out_5454),
            .b(out_21),
            .outp(out_5457)
        );        
        

        logic [WIDTH-1:0] out_5458;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5458 (
            .a(out_5456),
            .b(out_5457),
            .outp(out_5458)
        );        
        

        logic [WIDTH-1:0] out_5459;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.408)
        ) inst_5459 (
            .outp(out_5459)
        );
        

        logic [WIDTH-1:0] out_5460;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5460 (
            .a(out_3),
            .b(out_5459),
            .outp(out_5460)
        );        
        

        logic [WIDTH-1:0] out_5461;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5461 (
            .a(out_5458),
            .b(out_5460),
            .outp(out_5461)
        );        
        

        logic [WIDTH-1:0] out_5462;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5462 (
            .a(out_5461),
            .b(out_4559),
            .outp(out_5462)
        );        
        

        logic [WIDTH-1:0] out_5463;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5463 (
            .a(out_5462),
            .b(out_5447),
            .outp(out_5463)
        );        
        

        logic [WIDTH-1:0] out_5464;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5464 (
            .a(out_5449),
            .b(out_5463),
            .outp(out_5464)
        );        
        

        logic [WIDTH-1:0] out_5465;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.633)
        ) inst_5465 (
            .outp(out_5465)
        );
        

        logic [WIDTH-1:0] out_5466;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5466 (
            .a(out_5465),
            .b(out_3),
            .outp(out_5466)
        );        
        

        logic [WIDTH-1:0] out_5467;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5467 (
            .a(out_854),
            .b(out_5466),
            .outp(out_5467)
        );        
        

        logic [WIDTH-1:0] out_5468;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5468 (
            .a(out_5467),
            .b(out_4551),
            .outp(out_5468)
        );        
        

        logic [WIDTH-1:0] out_5469;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5469 (
            .a(out_5468),
            .b(out_4559),
            .outp(out_5469)
        );        
        

        logic [WIDTH-1:0] out_5470;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5470 (
            .a(out_5464),
            .b(out_5469),
            .outp(out_5470)
        );        
        

        logic [WIDTH-1:0] out_5471;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.1)
        ) inst_5471 (
            .outp(out_5471)
        );
        

        logic [WIDTH-1:0] out_5472;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5472 (
            .a(out_14),
            .b(out_5471),
            .outp(out_5472)
        );        
        

        logic [WIDTH-1:0] out_5473;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5473 (
            .in(out_5472),
            .outp(out_5473)
        );
        

        logic [WIDTH-1:0] out_5474;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.683)
        ) inst_5474 (
            .outp(out_5474)
        );
        

        logic [WIDTH-1:0] out_5475;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5475 (
            .a(out_3),
            .b(out_5474),
            .outp(out_5475)
        );        
        

        logic [WIDTH-1:0] out_5476;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5476 (
            .in(out_5475),
            .outp(out_5476)
        );
        

        logic [WIDTH-1:0] out_5477;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5477 (
            .a(out_5473),
            .b(out_5476),
            .outp(out_5477)
        );        
        

        logic [WIDTH-1:0] out_5478;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5478 (
            .in(out_5477),
            .outp(out_5478)
        );
        

        logic [WIDTH-1:0] out_5479;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5479 (
            .a(out_5478),
            .b(out_460),
            .outp(out_5479)
        );        
        

        logic [WIDTH-1:0] out_5480;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5480 (
            .a(out_5470),
            .b(out_5479),
            .outp(out_5480)
        );        
        

        logic [WIDTH-1:0] out_5481;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.75)
        ) inst_5481 (
            .outp(out_5481)
        );
        

        logic [WIDTH-1:0] out_5482;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5482 (
            .a(out_14),
            .b(out_5481),
            .outp(out_5482)
        );        
        

        logic [WIDTH-1:0] out_5483;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.508)
        ) inst_5483 (
            .outp(out_5483)
        );
        

        logic [WIDTH-1:0] out_5484;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5484 (
            .a(out_3),
            .b(out_5483),
            .outp(out_5484)
        );        
        

        logic [WIDTH-1:0] out_5485;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5485 (
            .a(out_5482),
            .b(out_5484),
            .outp(out_5485)
        );        
        

        logic [WIDTH-1:0] out_5486;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.408)
        ) inst_5486 (
            .outp(out_5486)
        );
        

        logic [WIDTH-1:0] out_5487;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5487 (
            .a(out_5486),
            .b(out_3),
            .outp(out_5487)
        );        
        

        logic [WIDTH-1:0] out_5488;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5488 (
            .a(out_5485),
            .b(out_5487),
            .outp(out_5488)
        );        
        

        logic [WIDTH-1:0] out_5489;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5489 (
            .a(out_5488),
            .b(out_4551),
            .outp(out_5489)
        );        
        

        logic [WIDTH-1:0] out_5490;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5490 (
            .a(out_5480),
            .b(out_5489),
            .outp(out_5490)
        );        
        

        logic [WIDTH-1:0] out_5491;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.258)
        ) inst_5491 (
            .outp(out_5491)
        );
        

        logic [WIDTH-1:0] out_5492;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5492 (
            .a(out_3),
            .b(out_5491),
            .outp(out_5492)
        );        
        

        logic [WIDTH-1:0] out_5493;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5493 (
            .a(out_5482),
            .b(out_5492),
            .outp(out_5493)
        );        
        

        logic [WIDTH-1:0] out_5494;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.158)
        ) inst_5494 (
            .outp(out_5494)
        );
        

        logic [WIDTH-1:0] out_5495;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5495 (
            .a(out_5494),
            .b(out_3),
            .outp(out_5495)
        );        
        

        logic [WIDTH-1:0] out_5496;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5496 (
            .a(out_5493),
            .b(out_5495),
            .outp(out_5496)
        );        
        

        logic [WIDTH-1:0] out_5497;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5497 (
            .a(out_5496),
            .b(out_4551),
            .outp(out_5497)
        );        
        

        logic [WIDTH-1:0] out_5498;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5498 (
            .a(out_5490),
            .b(out_5497),
            .outp(out_5498)
        );        
        

        logic [WIDTH-1:0] out_5499;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.925)
        ) inst_5499 (
            .outp(out_5499)
        );
        

        logic [WIDTH-1:0] out_5500;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5500 (
            .a(out_14),
            .b(out_5499),
            .outp(out_5500)
        );        
        

        logic [WIDTH-1:0] out_5501;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.008)
        ) inst_5501 (
            .outp(out_5501)
        );
        

        logic [WIDTH-1:0] out_5502;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5502 (
            .a(out_3),
            .b(out_5501),
            .outp(out_5502)
        );        
        

        logic [WIDTH-1:0] out_5503;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5503 (
            .a(out_5500),
            .b(out_5502),
            .outp(out_5503)
        );        
        

        logic [WIDTH-1:0] out_5504;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.908)
        ) inst_5504 (
            .outp(out_5504)
        );
        

        logic [WIDTH-1:0] out_5505;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5505 (
            .a(out_5504),
            .b(out_3),
            .outp(out_5505)
        );        
        

        logic [WIDTH-1:0] out_5506;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5506 (
            .a(out_5503),
            .b(out_5505),
            .outp(out_5506)
        );        
        

        logic [WIDTH-1:0] out_5507;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5507 (
            .a(out_5506),
            .b(out_4551),
            .outp(out_5507)
        );        
        

        logic [WIDTH-1:0] out_5508;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5508 (
            .a(out_5498),
            .b(out_5507),
            .outp(out_5508)
        );        
        

        logic [WIDTH-1:0] out_5509;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.05)
        ) inst_5509 (
            .outp(out_5509)
        );
        

        logic [WIDTH-1:0] out_5510;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5510 (
            .a(out_14),
            .b(out_5509),
            .outp(out_5510)
        );        
        

        logic [WIDTH-1:0] out_5511;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5511 (
            .a(out_5505),
            .b(out_5510),
            .outp(out_5511)
        );        
        

        logic [WIDTH-1:0] out_5512;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.75)
        ) inst_5512 (
            .outp(out_5512)
        );
        

        logic [WIDTH-1:0] out_5513;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5513 (
            .a(out_5512),
            .b(out_14),
            .outp(out_5513)
        );        
        

        logic [WIDTH-1:0] out_5514;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5514 (
            .a(out_5511),
            .b(out_5513),
            .outp(out_5514)
        );        
        

        logic [WIDTH-1:0] out_5515;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.558)
        ) inst_5515 (
            .outp(out_5515)
        );
        

        logic [WIDTH-1:0] out_5516;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5516 (
            .a(out_3),
            .b(out_5515),
            .outp(out_5516)
        );        
        

        logic [WIDTH-1:0] out_5517;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5517 (
            .a(out_5514),
            .b(out_5516),
            .outp(out_5517)
        );        
        

        logic [WIDTH-1:0] out_5518;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5518 (
            .in(out_5482),
            .outp(out_5518)
        );
        

        logic [WIDTH-1:0] out_5519;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.333)
        ) inst_5519 (
            .outp(out_5519)
        );
        

        logic [WIDTH-1:0] out_5520;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5520 (
            .a(out_3),
            .b(out_5519),
            .outp(out_5520)
        );        
        

        logic [WIDTH-1:0] out_5521;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5521 (
            .in(out_5520),
            .outp(out_5521)
        );
        

        logic [WIDTH-1:0] out_5522;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5522 (
            .a(out_5518),
            .b(out_5521),
            .outp(out_5522)
        );        
        

        logic [WIDTH-1:0] out_5523;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5523 (
            .in(out_5522),
            .outp(out_5523)
        );
        

        logic [WIDTH-1:0] out_5524;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5524 (
            .a(out_460),
            .b(out_5523),
            .outp(out_5524)
        );        
        

        logic [WIDTH-1:0] out_5525;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5525 (
            .a(out_5523),
            .b(out_9),
            .outp(out_5525)
        );        
        

        logic [WIDTH-1:0] out_5526;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5526 (
            .a(out_5524),
            .b(out_5525),
            .outp(out_5526)
        );        
        

        logic [WIDTH-1:0] out_5527;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.083)
        ) inst_5527 (
            .outp(out_5527)
        );
        

        logic [WIDTH-1:0] out_5528;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5528 (
            .a(out_3),
            .b(out_5527),
            .outp(out_5528)
        );        
        

        logic [WIDTH-1:0] out_5529;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5529 (
            .in(out_5528),
            .outp(out_5529)
        );
        

        logic [WIDTH-1:0] out_5530;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5530 (
            .a(out_5518),
            .b(out_5529),
            .outp(out_5530)
        );        
        

        logic [WIDTH-1:0] out_5531;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5531 (
            .in(out_5530),
            .outp(out_5531)
        );
        

        logic [WIDTH-1:0] out_5532;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5532 (
            .a(out_460),
            .b(out_5531),
            .outp(out_5532)
        );        
        

        logic [WIDTH-1:0] out_5533;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5533 (
            .a(out_5531),
            .b(out_9),
            .outp(out_5533)
        );        
        

        logic [WIDTH-1:0] out_5534;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5534 (
            .a(out_5532),
            .b(out_5533),
            .outp(out_5534)
        );        
        

        logic [WIDTH-1:0] out_5535;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5535 (
            .a(out_5526),
            .b(out_5534),
            .outp(out_5535)
        );        
        

        logic [WIDTH-1:0] out_5536;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5536 (
            .a(out_5517),
            .b(out_5535),
            .outp(out_5536)
        );        
        

        logic [WIDTH-1:0] out_5537;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5537 (
            .a(out_5508),
            .b(out_5536),
            .outp(out_5537)
        );        
        

        logic [WIDTH-1:0] out_5538;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5538 (
            .a(out_3044),
            .b(out_3384),
            .outp(out_5538)
        );        
        

        logic [WIDTH-1:0] out_5539;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5539 (
            .a(out_5538),
            .b(out_3582),
            .outp(out_5539)
        );        
        

        logic [WIDTH-1:0] out_5540;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5540 (
            .a(out_5539),
            .b(out_5350),
            .outp(out_5540)
        );        
        

        logic [WIDTH-1:0] out_5541;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.075)
        ) inst_5541 (
            .outp(out_5541)
        );
        

        logic [WIDTH-1:0] out_5542;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5542 (
            .a(out_5541),
            .b(out_3),
            .outp(out_5542)
        );        
        

        logic [WIDTH-1:0] out_5543;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5543 (
            .in(out_5542),
            .outp(out_5543)
        );
        

        logic [WIDTH-1:0] out_5544;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5544 (
            .a(out_3147),
            .b(out_5543),
            .outp(out_5544)
        );        
        

        logic [WIDTH-1:0] out_5545;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5545 (
            .in(out_5544),
            .outp(out_5545)
        );
        

        logic [WIDTH-1:0] out_5546;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5546 (
            .a(out_9),
            .b(out_5545),
            .outp(out_5546)
        );        
        

        logic [WIDTH-1:0] out_5547;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5547 (
            .a(out_5540),
            .b(out_5546),
            .outp(out_5547)
        );        
        

        logic [WIDTH-1:0] out_5548;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5548 (
            .a(out_5545),
            .b(out_21),
            .outp(out_5548)
        );        
        

        logic [WIDTH-1:0] out_5549;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5549 (
            .a(out_5547),
            .b(out_5548),
            .outp(out_5549)
        );        
        

        logic [WIDTH-1:0] out_5550;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5550 (
            .a(out_5537),
            .b(out_5549),
            .outp(out_5550)
        );        
        

        logic [WIDTH-1:0] out_5551;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5551 (
            .a(out_2782),
            .b(out_2786),
            .outp(out_5551)
        );        
        

        logic [WIDTH-1:0] out_5552;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5552 (
            .a(out_5551),
            .b(out_3297),
            .outp(out_5552)
        );        
        

        logic [WIDTH-1:0] out_5553;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5553 (
            .a(out_5552),
            .b(out_3299),
            .outp(out_5553)
        );        
        

        logic [WIDTH-1:0] out_5554;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5554 (
            .a(out_2790),
            .b(out_3147),
            .outp(out_5554)
        );        
        

        logic [WIDTH-1:0] out_5555;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5555 (
            .in(out_5554),
            .outp(out_5555)
        );
        

        logic [WIDTH-1:0] out_5556;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5556 (
            .a(out_5555),
            .b(out_21),
            .outp(out_5556)
        );        
        

        logic [WIDTH-1:0] out_5557;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.08)
        ) inst_5557 (
            .outp(out_5557)
        );
        

        logic [WIDTH-1:0] out_5558;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5558 (
            .a(out_5557),
            .b(out_556),
            .outp(out_5558)
        );        
        

        logic [WIDTH-1:0] out_5559;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5559 (
            .a(out_5558),
            .b(out_559),
            .outp(out_5559)
        );        
        

        logic [WIDTH-1:0] out_5560;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5560 (
            .a(out_3314),
            .b(out_5559),
            .outp(out_5560)
        );        
        

        logic [WIDTH-1:0] out_5561;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.885)
        ) inst_5561 (
            .outp(out_5561)
        );
        

        logic [WIDTH-1:0] out_5562;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5562 (
            .a(out_5561),
            .b(out_556),
            .outp(out_5562)
        );        
        

        logic [WIDTH-1:0] out_5563;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5563 (
            .a(out_5562),
            .b(out_566),
            .outp(out_5563)
        );        
        

        logic [WIDTH-1:0] out_5564;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5564 (
            .in(out_5563),
            .outp(out_5564)
        );
        

        logic [WIDTH-1:0] out_5565;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5565 (
            .a(out_5560),
            .b(out_5564),
            .outp(out_5565)
        );        
        

        logic [WIDTH-1:0] out_5566;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.885)
        ) inst_5566 (
            .outp(out_5566)
        );
        

        logic [WIDTH-1:0] out_5567;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5567 (
            .a(out_5566),
            .b(out_556),
            .outp(out_5567)
        );        
        

        logic [WIDTH-1:0] out_5568;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5568 (
            .a(out_5567),
            .b(out_566),
            .outp(out_5568)
        );        
        

        logic [WIDTH-1:0] out_5569;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5569 (
            .a(out_3325),
            .b(out_5568),
            .outp(out_5569)
        );        
        

        logic [WIDTH-1:0] out_5570;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.08)
        ) inst_5570 (
            .outp(out_5570)
        );
        

        logic [WIDTH-1:0] out_5571;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5571 (
            .a(out_5570),
            .b(out_556),
            .outp(out_5571)
        );        
        

        logic [WIDTH-1:0] out_5572;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5572 (
            .a(out_559),
            .b(out_5571),
            .outp(out_5572)
        );        
        

        logic [WIDTH-1:0] out_5573;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5573 (
            .a(out_5569),
            .b(out_5572),
            .outp(out_5573)
        );        
        

        logic [WIDTH-1:0] out_5574;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5574 (
            .a(out_5565),
            .b(out_5573),
            .outp(out_5574)
        );        
        

        logic [WIDTH-1:0] out_5575;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5575 (
            .in(out_5574),
            .outp(out_5575)
        );
        

        logic [WIDTH-1:0] out_5576;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5576 (
            .a(out_5556),
            .b(out_5575),
            .outp(out_5576)
        );        
        

        logic [WIDTH-1:0] out_5577;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5577 (
            .a(out_9),
            .b(out_5555),
            .outp(out_5577)
        );        
        

        logic [WIDTH-1:0] out_5578;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5578 (
            .a(out_5576),
            .b(out_5577),
            .outp(out_5578)
        );        
        

        logic [WIDTH-1:0] out_5579;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5579 (
            .a(out_5553),
            .b(out_5578),
            .outp(out_5579)
        );        
        

        logic [WIDTH-1:0] out_5580;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5580 (
            .a(out_5556),
            .b(out_5579),
            .outp(out_5580)
        );        
        

        logic [WIDTH-1:0] out_5581;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5581 (
            .a(out_5550),
            .b(out_5580),
            .outp(out_5581)
        );        
        

        logic [WIDTH-1:0] out_5582;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.715)
        ) inst_5582 (
            .outp(out_5582)
        );
        

        logic [WIDTH-1:0] out_5583;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5583 (
            .a(out_14),
            .b(out_5582),
            .outp(out_5583)
        );        
        

        logic [WIDTH-1:0] out_5584;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.625)
        ) inst_5584 (
            .outp(out_5584)
        );
        

        logic [WIDTH-1:0] out_5585;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5585 (
            .a(out_5584),
            .b(out_14),
            .outp(out_5585)
        );        
        

        logic [WIDTH-1:0] out_5586;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5586 (
            .a(out_5583),
            .b(out_5585),
            .outp(out_5586)
        );        
        

        logic [WIDTH-1:0] out_5587;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.058)
        ) inst_5587 (
            .outp(out_5587)
        );
        

        logic [WIDTH-1:0] out_5588;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5588 (
            .a(out_3),
            .b(out_5587),
            .outp(out_5588)
        );        
        

        logic [WIDTH-1:0] out_5589;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5589 (
            .a(out_5586),
            .b(out_5588),
            .outp(out_5589)
        );        
        

        logic [WIDTH-1:0] out_5590;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.558)
        ) inst_5590 (
            .outp(out_5590)
        );
        

        logic [WIDTH-1:0] out_5591;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5591 (
            .a(out_5590),
            .b(out_3),
            .outp(out_5591)
        );        
        

        logic [WIDTH-1:0] out_5592;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5592 (
            .a(out_5589),
            .b(out_5591),
            .outp(out_5592)
        );        
        

        logic [WIDTH-1:0] out_5593;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.783)
        ) inst_5593 (
            .outp(out_5593)
        );
        

        logic [WIDTH-1:0] out_5594;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5594 (
            .a(out_3),
            .b(out_5593),
            .outp(out_5594)
        );        
        

        logic [WIDTH-1:0] out_5595;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5595 (
            .in(out_5594),
            .outp(out_5595)
        );
        

        logic [WIDTH-1:0] out_5596;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5596 (
            .a(out_4534),
            .b(out_5595),
            .outp(out_5596)
        );        
        

        logic [WIDTH-1:0] out_5597;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5597 (
            .in(out_5596),
            .outp(out_5597)
        );
        

        logic [WIDTH-1:0] out_5598;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5598 (
            .a(out_5597),
            .b(out_21),
            .outp(out_5598)
        );        
        

        logic [WIDTH-1:0] out_5599;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.08875)
        ) inst_5599 (
            .outp(out_5599)
        );
        

        logic [WIDTH-1:0] out_5600;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5600 (
            .a(out_553),
            .b(out_5599),
            .outp(out_5600)
        );        
        

        logic [WIDTH-1:0] out_5601;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.7447)
        ) inst_5601 (
            .outp(out_5601)
        );
        

        logic [WIDTH-1:0] out_5602;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5602 (
            .a(out_559),
            .b(out_5601),
            .outp(out_5602)
        );        
        

        logic [WIDTH-1:0] out_5603;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5603 (
            .a(out_556),
            .b(out_5602),
            .outp(out_5603)
        );        
        

        logic [WIDTH-1:0] out_5604;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5604 (
            .a(out_5600),
            .b(out_5603),
            .outp(out_5604)
        );        
        

        logic [WIDTH-1:0] out_5605;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6547)
        ) inst_5605 (
            .outp(out_5605)
        );
        

        logic [WIDTH-1:0] out_5606;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5606 (
            .a(out_5605),
            .b(out_2653),
            .outp(out_5606)
        );        
        

        logic [WIDTH-1:0] out_5607;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5607 (
            .a(out_5604),
            .b(out_5606),
            .outp(out_5607)
        );        
        

        logic [WIDTH-1:0] out_5608;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5608 (
            .a(out_2653),
            .b(out_5605),
            .outp(out_5608)
        );        
        

        logic [WIDTH-1:0] out_5609;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5609 (
            .a(out_5602),
            .b(out_556),
            .outp(out_5609)
        );        
        

        logic [WIDTH-1:0] out_5610;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5610 (
            .a(out_5608),
            .b(out_5609),
            .outp(out_5610)
        );        
        

        logic [WIDTH-1:0] out_5611;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5611 (
            .a(out_5599),
            .b(out_553),
            .outp(out_5611)
        );        
        

        logic [WIDTH-1:0] out_5612;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5612 (
            .a(out_5610),
            .b(out_5611),
            .outp(out_5612)
        );        
        

        logic [WIDTH-1:0] out_5613;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5613 (
            .a(out_5607),
            .b(out_5612),
            .outp(out_5613)
        );        
        

        logic [WIDTH-1:0] out_5614;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5614 (
            .in(out_5613),
            .outp(out_5614)
        );
        

        logic [WIDTH-1:0] out_5615;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5615 (
            .a(out_5598),
            .b(out_5614),
            .outp(out_5615)
        );        
        

        logic [WIDTH-1:0] out_5616;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5616 (
            .a(out_9),
            .b(out_5597),
            .outp(out_5616)
        );        
        

        logic [WIDTH-1:0] out_5617;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5617 (
            .a(out_5615),
            .b(out_5616),
            .outp(out_5617)
        );        
        

        logic [WIDTH-1:0] out_5618;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5618 (
            .a(out_5592),
            .b(out_5617),
            .outp(out_5618)
        );        
        

        logic [WIDTH-1:0] out_5619;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5619 (
            .a(out_5598),
            .b(out_5618),
            .outp(out_5619)
        );        
        

        logic [WIDTH-1:0] out_5620;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5620 (
            .a(out_5581),
            .b(out_5619),
            .outp(out_5620)
        );        
        

        logic [WIDTH-1:0] out_5621;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5621 (
            .a(out_4548),
            .b(out_4551),
            .outp(out_5621)
        );        
        

        logic [WIDTH-1:0] out_5622;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5622 (
            .a(out_5621),
            .b(out_5460),
            .outp(out_5622)
        );        
        

        logic [WIDTH-1:0] out_5623;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.308)
        ) inst_5623 (
            .outp(out_5623)
        );
        

        logic [WIDTH-1:0] out_5624;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5624 (
            .a(out_5623),
            .b(out_3),
            .outp(out_5624)
        );        
        

        logic [WIDTH-1:0] out_5625;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5625 (
            .a(out_5622),
            .b(out_5624),
            .outp(out_5625)
        );        
        

        logic [WIDTH-1:0] out_5626;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5626 (
            .a(out_5620),
            .b(out_5625),
            .outp(out_5626)
        );        
        

        logic [WIDTH-1:0] out_5627;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5627 (
            .a(out_3),
            .b(out_220),
            .outp(out_5627)
        );        
        

        logic [WIDTH-1:0] out_5628;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5628 (
            .in(out_5627),
            .outp(out_5628)
        );
        

        logic [WIDTH-1:0] out_5629;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5629 (
            .a(out_4534),
            .b(out_5628),
            .outp(out_5629)
        );        
        

        logic [WIDTH-1:0] out_5630;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5630 (
            .in(out_5629),
            .outp(out_5630)
        );
        

        logic [WIDTH-1:0] out_5631;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5631 (
            .a(out_5630),
            .b(out_21),
            .outp(out_5631)
        );        
        

        logic [WIDTH-1:0] out_5632;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5632 (
            .a(out_9),
            .b(out_5630),
            .outp(out_5632)
        );        
        

        logic [WIDTH-1:0] out_5633;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5633 (
            .a(out_5631),
            .b(out_5632),
            .outp(out_5633)
        );        
        

        logic [WIDTH-1:0] out_5634;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5634 (
            .a(out_5626),
            .b(out_5633),
            .outp(out_5634)
        );        
        

        logic [WIDTH-1:0] out_5635;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.8325)
        ) inst_5635 (
            .outp(out_5635)
        );
        

        logic [WIDTH-1:0] out_5636;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5636 (
            .a(out_5635),
            .b(out_131),
            .outp(out_5636)
        );        
        

        logic [WIDTH-1:0] out_5637;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5637 (
            .a(out_127),
            .b(out_5636),
            .outp(out_5637)
        );        
        

        logic [WIDTH-1:0] out_5638;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5638 (
            .a(out_4508),
            .b(out_5637),
            .outp(out_5638)
        );        
        

        logic [WIDTH-1:0] out_5639;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6375)
        ) inst_5639 (
            .outp(out_5639)
        );
        

        logic [WIDTH-1:0] out_5640;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5640 (
            .a(out_5639),
            .b(out_124),
            .outp(out_5640)
        );        
        

        logic [WIDTH-1:0] out_5641;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5641 (
            .a(out_5640),
            .b(out_127),
            .outp(out_5641)
        );        
        

        logic [WIDTH-1:0] out_5642;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5642 (
            .a(out_5638),
            .b(out_5641),
            .outp(out_5642)
        );        
        

        logic [WIDTH-1:0] out_5643;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5643 (
            .a(out_5634),
            .b(out_5642),
            .outp(out_5643)
        );        
        

        logic [WIDTH-1:0] out_5644;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5644 (
            .a(out_127),
            .b(out_5640),
            .outp(out_5644)
        );        
        

        logic [WIDTH-1:0] out_5645;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5645 (
            .a(out_5636),
            .b(out_127),
            .outp(out_5645)
        );        
        

        logic [WIDTH-1:0] out_5646;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5646 (
            .a(out_5644),
            .b(out_5645),
            .outp(out_5646)
        );        
        

        logic [WIDTH-1:0] out_5647;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5647 (
            .a(out_5646),
            .b(out_4513),
            .outp(out_5647)
        );        
        

        logic [WIDTH-1:0] out_5648;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5648 (
            .a(out_5643),
            .b(out_5647),
            .outp(out_5648)
        );        
        

        logic [WIDTH-1:0] out_5649;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5649 (
            .a(out_5644),
            .b(out_4521),
            .outp(out_5649)
        );        
        

        logic [WIDTH-1:0] out_5650;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.7775)
        ) inst_5650 (
            .outp(out_5650)
        );
        

        logic [WIDTH-1:0] out_5651;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5651 (
            .a(out_5650),
            .b(out_131),
            .outp(out_5651)
        );        
        

        logic [WIDTH-1:0] out_5652;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5652 (
            .a(out_5651),
            .b(out_127),
            .outp(out_5652)
        );        
        

        logic [WIDTH-1:0] out_5653;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5653 (
            .a(out_5649),
            .b(out_5652),
            .outp(out_5653)
        );        
        

        logic [WIDTH-1:0] out_5654;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5654 (
            .a(out_5648),
            .b(out_5653),
            .outp(out_5654)
        );        
        

        logic [WIDTH-1:0] out_5655;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5655 (
            .a(out_127),
            .b(out_5651),
            .outp(out_5655)
        );        
        

        logic [WIDTH-1:0] out_5656;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5656 (
            .a(out_5641),
            .b(out_5655),
            .outp(out_5656)
        );        
        

        logic [WIDTH-1:0] out_5657;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5657 (
            .a(out_5656),
            .b(out_4526),
            .outp(out_5657)
        );        
        

        logic [WIDTH-1:0] out_5658;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5658 (
            .a(out_5654),
            .b(out_5657),
            .outp(out_5658)
        );        
        

        logic [WIDTH-1:0] out_5659;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.4775)
        ) inst_5659 (
            .outp(out_5659)
        );
        

        logic [WIDTH-1:0] out_5660;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5660 (
            .a(out_5659),
            .b(out_4477),
            .outp(out_5660)
        );        
        

        logic [WIDTH-1:0] out_5661;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5661 (
            .a(out_4508),
            .b(out_5660),
            .outp(out_5661)
        );        
        

        logic [WIDTH-1:0] out_5662;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.6725)
        ) inst_5662 (
            .outp(out_5662)
        );
        

        logic [WIDTH-1:0] out_5663;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5663 (
            .a(out_4480),
            .b(out_5662),
            .outp(out_5663)
        );        
        

        logic [WIDTH-1:0] out_5664;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5664 (
            .a(out_5661),
            .b(out_5663),
            .outp(out_5664)
        );        
        

        logic [WIDTH-1:0] out_5665;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5665 (
            .a(out_5658),
            .b(out_5664),
            .outp(out_5665)
        );        
        

        logic [WIDTH-1:0] out_5666;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5666 (
            .a(out_5662),
            .b(out_4480),
            .outp(out_5666)
        );        
        

        logic [WIDTH-1:0] out_5667;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5667 (
            .a(out_4513),
            .b(out_5666),
            .outp(out_5667)
        );        
        

        logic [WIDTH-1:0] out_5668;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5668 (
            .a(out_4477),
            .b(out_5659),
            .outp(out_5668)
        );        
        

        logic [WIDTH-1:0] out_5669;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5669 (
            .a(out_5667),
            .b(out_5668),
            .outp(out_5669)
        );        
        

        logic [WIDTH-1:0] out_5670;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5670 (
            .a(out_5665),
            .b(out_5669),
            .outp(out_5670)
        );        
        

        logic [WIDTH-1:0] out_5671;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5671 (
            .a(out_4521),
            .b(out_5666),
            .outp(out_5671)
        );        
        

        logic [WIDTH-1:0] out_5672;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5325)
        ) inst_5672 (
            .outp(out_5672)
        );
        

        logic [WIDTH-1:0] out_5673;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5673 (
            .a(out_4477),
            .b(out_5672),
            .outp(out_5673)
        );        
        

        logic [WIDTH-1:0] out_5674;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5674 (
            .a(out_5671),
            .b(out_5673),
            .outp(out_5674)
        );        
        

        logic [WIDTH-1:0] out_5675;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5675 (
            .a(out_5670),
            .b(out_5674),
            .outp(out_5675)
        );        
        

        logic [WIDTH-1:0] out_5676;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5676 (
            .a(out_4526),
            .b(out_5663),
            .outp(out_5676)
        );        
        

        logic [WIDTH-1:0] out_5677;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5677 (
            .a(out_5672),
            .b(out_4477),
            .outp(out_5677)
        );        
        

        logic [WIDTH-1:0] out_5678;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5678 (
            .a(out_5676),
            .b(out_5677),
            .outp(out_5678)
        );        
        

        logic [WIDTH-1:0] out_5679;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5679 (
            .a(out_5675),
            .b(out_5678),
            .outp(out_5679)
        );        
        

        logic [WIDTH-1:0] out_5680;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5575)
        ) inst_5680 (
            .outp(out_5680)
        );
        

        logic [WIDTH-1:0] out_5681;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5681 (
            .a(out_5680),
            .b(out_131),
            .outp(out_5681)
        );        
        

        logic [WIDTH-1:0] out_5682;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5682 (
            .a(out_127),
            .b(out_5681),
            .outp(out_5682)
        );        
        

        logic [WIDTH-1:0] out_5683;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5683 (
            .a(out_4508),
            .b(out_5682),
            .outp(out_5683)
        );        
        

        logic [WIDTH-1:0] out_5684;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.3625)
        ) inst_5684 (
            .outp(out_5684)
        );
        

        logic [WIDTH-1:0] out_5685;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5685 (
            .a(out_5684),
            .b(out_124),
            .outp(out_5685)
        );        
        

        logic [WIDTH-1:0] out_5686;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5686 (
            .a(out_5685),
            .b(out_127),
            .outp(out_5686)
        );        
        

        logic [WIDTH-1:0] out_5687;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5687 (
            .a(out_5683),
            .b(out_5686),
            .outp(out_5687)
        );        
        

        logic [WIDTH-1:0] out_5688;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5688 (
            .a(out_5679),
            .b(out_5687),
            .outp(out_5688)
        );        
        

        logic [WIDTH-1:0] out_5689;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5689 (
            .a(out_127),
            .b(out_5685),
            .outp(out_5689)
        );        
        

        logic [WIDTH-1:0] out_5690;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5690 (
            .a(out_4513),
            .b(out_5689),
            .outp(out_5690)
        );        
        

        logic [WIDTH-1:0] out_5691;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5691 (
            .a(out_5681),
            .b(out_127),
            .outp(out_5691)
        );        
        

        logic [WIDTH-1:0] out_5692;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5692 (
            .a(out_5690),
            .b(out_5691),
            .outp(out_5692)
        );        
        

        logic [WIDTH-1:0] out_5693;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5693 (
            .a(out_5688),
            .b(out_5692),
            .outp(out_5693)
        );        
        

        logic [WIDTH-1:0] out_5694;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5694 (
            .a(out_4521),
            .b(out_5689),
            .outp(out_5694)
        );        
        

        logic [WIDTH-1:0] out_5695;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5025)
        ) inst_5695 (
            .outp(out_5695)
        );
        

        logic [WIDTH-1:0] out_5696;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5696 (
            .a(out_5695),
            .b(out_131),
            .outp(out_5696)
        );        
        

        logic [WIDTH-1:0] out_5697;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5697 (
            .a(out_5696),
            .b(out_127),
            .outp(out_5697)
        );        
        

        logic [WIDTH-1:0] out_5698;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5698 (
            .a(out_5694),
            .b(out_5697),
            .outp(out_5698)
        );        
        

        logic [WIDTH-1:0] out_5699;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5699 (
            .a(out_5693),
            .b(out_5698),
            .outp(out_5699)
        );        
        

        logic [WIDTH-1:0] out_5700;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5700 (
            .a(out_4526),
            .b(out_5686),
            .outp(out_5700)
        );        
        

        logic [WIDTH-1:0] out_5701;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5701 (
            .a(out_127),
            .b(out_5696),
            .outp(out_5701)
        );        
        

        logic [WIDTH-1:0] out_5702;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5702 (
            .a(out_5700),
            .b(out_5701),
            .outp(out_5702)
        );        
        

        logic [WIDTH-1:0] out_5703;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5703 (
            .a(out_5699),
            .b(out_5702),
            .outp(out_5703)
        );        
        

        logic [WIDTH-1:0] out_5704;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2025)
        ) inst_5704 (
            .outp(out_5704)
        );
        

        logic [WIDTH-1:0] out_5705;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5705 (
            .a(out_5704),
            .b(out_4477),
            .outp(out_5705)
        );        
        

        logic [WIDTH-1:0] out_5706;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5706 (
            .a(out_4508),
            .b(out_5705),
            .outp(out_5706)
        );        
        

        logic [WIDTH-1:0] out_5707;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.3975)
        ) inst_5707 (
            .outp(out_5707)
        );
        

        logic [WIDTH-1:0] out_5708;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5708 (
            .a(out_4480),
            .b(out_5707),
            .outp(out_5708)
        );        
        

        logic [WIDTH-1:0] out_5709;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5709 (
            .a(out_5706),
            .b(out_5708),
            .outp(out_5709)
        );        
        

        logic [WIDTH-1:0] out_5710;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5710 (
            .a(out_5703),
            .b(out_5709),
            .outp(out_5710)
        );        
        

        logic [WIDTH-1:0] out_5711;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5711 (
            .a(out_5707),
            .b(out_4480),
            .outp(out_5711)
        );        
        

        logic [WIDTH-1:0] out_5712;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5712 (
            .a(out_4513),
            .b(out_5711),
            .outp(out_5712)
        );        
        

        logic [WIDTH-1:0] out_5713;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5713 (
            .a(out_4477),
            .b(out_5704),
            .outp(out_5713)
        );        
        

        logic [WIDTH-1:0] out_5714;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5714 (
            .a(out_5712),
            .b(out_5713),
            .outp(out_5714)
        );        
        

        logic [WIDTH-1:0] out_5715;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5715 (
            .a(out_5710),
            .b(out_5714),
            .outp(out_5715)
        );        
        

        logic [WIDTH-1:0] out_5716;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5716 (
            .a(out_4521),
            .b(out_5711),
            .outp(out_5716)
        );        
        

        logic [WIDTH-1:0] out_5717;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2575)
        ) inst_5717 (
            .outp(out_5717)
        );
        

        logic [WIDTH-1:0] out_5718;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5718 (
            .a(out_4477),
            .b(out_5717),
            .outp(out_5718)
        );        
        

        logic [WIDTH-1:0] out_5719;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5719 (
            .a(out_5716),
            .b(out_5718),
            .outp(out_5719)
        );        
        

        logic [WIDTH-1:0] out_5720;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5720 (
            .a(out_5715),
            .b(out_5719),
            .outp(out_5720)
        );        
        

        logic [WIDTH-1:0] out_5721;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5721 (
            .a(out_4526),
            .b(out_5708),
            .outp(out_5721)
        );        
        

        logic [WIDTH-1:0] out_5722;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5722 (
            .a(out_5717),
            .b(out_4477),
            .outp(out_5722)
        );        
        

        logic [WIDTH-1:0] out_5723;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5723 (
            .a(out_5721),
            .b(out_5722),
            .outp(out_5723)
        );        
        

        logic [WIDTH-1:0] out_5724;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5724 (
            .a(out_5720),
            .b(out_5723),
            .outp(out_5724)
        );        
        

        logic [WIDTH-1:0] out_5725;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.224999)
        ) inst_5725 (
            .outp(out_5725)
        );
        

        logic [WIDTH-1:0] out_5726;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5726 (
            .a(out_3),
            .b(out_5725),
            .outp(out_5726)
        );        
        

        logic [WIDTH-1:0] out_5727;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5727 (
            .in(out_5726),
            .outp(out_5727)
        );
        

        logic [WIDTH-1:0] out_5728;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5728 (
            .a(out_4534),
            .b(out_5727),
            .outp(out_5728)
        );        
        

        logic [WIDTH-1:0] out_5729;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5729 (
            .in(out_5728),
            .outp(out_5729)
        );
        

        logic [WIDTH-1:0] out_5730;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5730 (
            .a(out_9),
            .b(out_5729),
            .outp(out_5730)
        );        
        

        logic [WIDTH-1:0] out_5731;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5731 (
            .a(out_5729),
            .b(out_21),
            .outp(out_5731)
        );        
        

        logic [WIDTH-1:0] out_5732;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5732 (
            .a(out_5730),
            .b(out_5731),
            .outp(out_5732)
        );        
        

        logic [WIDTH-1:0] out_5733;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5733 (
            .a(out_5724),
            .b(out_5732),
            .outp(out_5733)
        );        
        

        logic [WIDTH-1:0] out_5734;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2)
        ) inst_5734 (
            .outp(out_5734)
        );
        

        logic [WIDTH-1:0] out_5735;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5735 (
            .a(out_566),
            .b(out_5734),
            .outp(out_5735)
        );        
        

        logic [WIDTH-1:0] out_5736;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.104)
        ) inst_5736 (
            .outp(out_5736)
        );
        

        logic [WIDTH-1:0] out_5737;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5737 (
            .a(out_862),
            .b(out_5736),
            .outp(out_5737)
        );        
        

        logic [WIDTH-1:0] out_5738;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5738 (
            .a(out_5735),
            .b(out_5737),
            .outp(out_5738)
        );        
        

        logic [WIDTH-1:0] out_5739;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.054)
        ) inst_5739 (
            .outp(out_5739)
        );
        

        logic [WIDTH-1:0] out_5740;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5740 (
            .a(out_5739),
            .b(out_868),
            .outp(out_5740)
        );        
        

        logic [WIDTH-1:0] out_5741;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5741 (
            .a(out_5738),
            .b(out_5740),
            .outp(out_5741)
        );        
        

        logic [WIDTH-1:0] out_5742;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5742 (
            .a(out_868),
            .b(out_5739),
            .outp(out_5742)
        );        
        

        logic [WIDTH-1:0] out_5743;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5743 (
            .a(out_5736),
            .b(out_862),
            .outp(out_5743)
        );        
        

        logic [WIDTH-1:0] out_5744;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5744 (
            .a(out_5742),
            .b(out_5743),
            .outp(out_5744)
        );        
        

        logic [WIDTH-1:0] out_5745;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5745 (
            .a(out_5734),
            .b(out_566),
            .outp(out_5745)
        );        
        

        logic [WIDTH-1:0] out_5746;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5746 (
            .a(out_5744),
            .b(out_5745),
            .outp(out_5746)
        );        
        

        logic [WIDTH-1:0] out_5747;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5747 (
            .a(out_5741),
            .b(out_5746),
            .outp(out_5747)
        );        
        

        logic [WIDTH-1:0] out_5748;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.968)
        ) inst_5748 (
            .outp(out_5748)
        );
        

        logic [WIDTH-1:0] out_5749;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5749 (
            .a(out_878),
            .b(out_5748),
            .outp(out_5749)
        );        
        

        logic [WIDTH-1:0] out_5750;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5750 (
            .a(out_3),
            .b(out_5749),
            .outp(out_5750)
        );        
        

        logic [WIDTH-1:0] out_5751;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.8858)
        ) inst_5751 (
            .outp(out_5751)
        );
        

        logic [WIDTH-1:0] out_5752;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5752 (
            .a(out_884),
            .b(out_886),
            .outp(out_5752)
        );        
        

        logic [WIDTH-1:0] out_5753;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5753 (
            .a(out_5751),
            .b(out_5752),
            .outp(out_5753)
        );        
        

        logic [WIDTH-1:0] out_5754;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5754 (
            .a(out_5750),
            .b(out_5753),
            .outp(out_5754)
        );        
        

        logic [WIDTH-1:0] out_5755;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.7272)
        ) inst_5755 (
            .outp(out_5755)
        );
        

        logic [WIDTH-1:0] out_5756;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5756 (
            .a(out_5755),
            .b(out_891),
            .outp(out_5756)
        );        
        

        logic [WIDTH-1:0] out_5757;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5757 (
            .a(out_5756),
            .b(out_894),
            .outp(out_5757)
        );        
        

        logic [WIDTH-1:0] out_5758;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5758 (
            .a(out_5754),
            .b(out_5757),
            .outp(out_5758)
        );        
        

        logic [WIDTH-1:0] out_5759;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5759 (
            .a(out_5747),
            .b(out_5758),
            .outp(out_5759)
        );        
        

        logic [WIDTH-1:0] out_5760;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5760 (
            .a(out_894),
            .b(out_5756),
            .outp(out_5760)
        );        
        

        logic [WIDTH-1:0] out_5761;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5761 (
            .a(out_5752),
            .b(out_5751),
            .outp(out_5761)
        );        
        

        logic [WIDTH-1:0] out_5762;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5762 (
            .a(out_5760),
            .b(out_5761),
            .outp(out_5762)
        );        
        

        logic [WIDTH-1:0] out_5763;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5763 (
            .a(out_5749),
            .b(out_3),
            .outp(out_5763)
        );        
        

        logic [WIDTH-1:0] out_5764;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5764 (
            .a(out_5762),
            .b(out_5763),
            .outp(out_5764)
        );        
        

        logic [WIDTH-1:0] out_5765;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5765 (
            .a(out_5759),
            .b(out_5764),
            .outp(out_5765)
        );        
        

        logic [WIDTH-1:0] out_5766;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.351)
        ) inst_5766 (
            .outp(out_5766)
        );
        

        logic [WIDTH-1:0] out_5767;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5767 (
            .a(out_5766),
            .b(out_910),
            .outp(out_5767)
        );        
        

        logic [WIDTH-1:0] out_5768;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2978)
        ) inst_5768 (
            .outp(out_5768)
        );
        

        logic [WIDTH-1:0] out_5769;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5769 (
            .a(out_5768),
            .b(out_886),
            .outp(out_5769)
        );        
        

        logic [WIDTH-1:0] out_5770;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5770 (
            .a(out_5767),
            .b(out_5769),
            .outp(out_5770)
        );        
        

        logic [WIDTH-1:0] out_5771;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.7433)
        ) inst_5771 (
            .outp(out_5771)
        );
        

        logic [WIDTH-1:0] out_5772;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5772 (
            .a(out_916),
            .b(out_5771),
            .outp(out_5772)
        );        
        

        logic [WIDTH-1:0] out_5773;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5773 (
            .a(out_5770),
            .b(out_5772),
            .outp(out_5773)
        );        
        

        logic [WIDTH-1:0] out_5774;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5774 (
            .a(out_5765),
            .b(out_5773),
            .outp(out_5774)
        );        
        

        logic [WIDTH-1:0] out_5775;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5775 (
            .a(out_5771),
            .b(out_916),
            .outp(out_5775)
        );        
        

        logic [WIDTH-1:0] out_5776;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5776 (
            .a(out_886),
            .b(out_5768),
            .outp(out_5776)
        );        
        

        logic [WIDTH-1:0] out_5777;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5777 (
            .a(out_5775),
            .b(out_5776),
            .outp(out_5777)
        );        
        

        logic [WIDTH-1:0] out_5778;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5778 (
            .a(out_910),
            .b(out_5766),
            .outp(out_5778)
        );        
        

        logic [WIDTH-1:0] out_5779;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5779 (
            .a(out_5777),
            .b(out_5778),
            .outp(out_5779)
        );        
        

        logic [WIDTH-1:0] out_5780;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5780 (
            .a(out_5774),
            .b(out_5779),
            .outp(out_5780)
        );        
        

        logic [WIDTH-1:0] out_5781;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.96)
        ) inst_5781 (
            .outp(out_5781)
        );
        

        logic [WIDTH-1:0] out_5782;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5782 (
            .a(out_928),
            .b(out_5781),
            .outp(out_5782)
        );        
        

        logic [WIDTH-1:0] out_5783;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2994)
        ) inst_5783 (
            .outp(out_5783)
        );
        

        logic [WIDTH-1:0] out_5784;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5784 (
            .a(out_5783),
            .b(out_928),
            .outp(out_5784)
        );        
        

        logic [WIDTH-1:0] out_5785;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5785 (
            .a(out_127),
            .b(out_5784),
            .outp(out_5785)
        );        
        

        logic [WIDTH-1:0] out_5786;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5786 (
            .a(out_5782),
            .b(out_5785),
            .outp(out_5786)
        );        
        

        logic [WIDTH-1:0] out_5787;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.0394)
        ) inst_5787 (
            .outp(out_5787)
        );
        

        logic [WIDTH-1:0] out_5788;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5788 (
            .a(out_5787),
            .b(out_127),
            .outp(out_5788)
        );        
        

        logic [WIDTH-1:0] out_5789;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5789 (
            .a(out_5786),
            .b(out_5788),
            .outp(out_5789)
        );        
        

        logic [WIDTH-1:0] out_5790;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5790 (
            .a(out_5780),
            .b(out_5789),
            .outp(out_5790)
        );        
        

        logic [WIDTH-1:0] out_5791;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5791 (
            .a(out_127),
            .b(out_5787),
            .outp(out_5791)
        );        
        

        logic [WIDTH-1:0] out_5792;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5792 (
            .a(out_5784),
            .b(out_127),
            .outp(out_5792)
        );        
        

        logic [WIDTH-1:0] out_5793;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5793 (
            .a(out_5791),
            .b(out_5792),
            .outp(out_5793)
        );        
        

        logic [WIDTH-1:0] out_5794;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5794 (
            .a(out_5781),
            .b(out_928),
            .outp(out_5794)
        );        
        

        logic [WIDTH-1:0] out_5795;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5795 (
            .a(out_5793),
            .b(out_5794),
            .outp(out_5795)
        );        
        

        logic [WIDTH-1:0] out_5796;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5796 (
            .a(out_5790),
            .b(out_5795),
            .outp(out_5796)
        );        
        

        logic [WIDTH-1:0] out_5797;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5797 (
            .in(out_5796),
            .outp(out_5797)
        );
        

        logic [WIDTH-1:0] out_5798;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5798 (
            .a(out_4551),
            .b(out_5797),
            .outp(out_5798)
        );        
        

        logic [WIDTH-1:0] out_5799;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.4)
        ) inst_5799 (
            .outp(out_5799)
        );
        

        logic [WIDTH-1:0] out_5800;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5800 (
            .a(out_14),
            .b(out_5799),
            .outp(out_5800)
        );        
        

        logic [WIDTH-1:0] out_5801;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5801 (
            .a(out_5798),
            .b(out_5800),
            .outp(out_5801)
        );        
        

        logic [WIDTH-1:0] out_5802;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.108)
        ) inst_5802 (
            .outp(out_5802)
        );
        

        logic [WIDTH-1:0] out_5803;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5803 (
            .a(out_3),
            .b(out_5802),
            .outp(out_5803)
        );        
        

        logic [WIDTH-1:0] out_5804;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5804 (
            .a(out_5801),
            .b(out_5803),
            .outp(out_5804)
        );        
        

        logic [WIDTH-1:0] out_5805;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.608)
        ) inst_5805 (
            .outp(out_5805)
        );
        

        logic [WIDTH-1:0] out_5806;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5806 (
            .a(out_5805),
            .b(out_3),
            .outp(out_5806)
        );        
        

        logic [WIDTH-1:0] out_5807;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5807 (
            .a(out_5804),
            .b(out_5806),
            .outp(out_5807)
        );        
        

        logic [WIDTH-1:0] out_5808;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5808 (
            .a(out_5733),
            .b(out_5807),
            .outp(out_5808)
        );        
        

        logic [WIDTH-1:0] out_5809;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.25)
        ) inst_5809 (
            .outp(out_5809)
        );
        

        logic [WIDTH-1:0] out_5810;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5810 (
            .a(out_3),
            .b(out_5809),
            .outp(out_5810)
        );        
        

        logic [WIDTH-1:0] out_5811;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5811 (
            .a(out_5442),
            .b(out_5810),
            .outp(out_5811)
        );        
        

        logic [WIDTH-1:0] out_5812;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.15)
        ) inst_5812 (
            .outp(out_5812)
        );
        

        logic [WIDTH-1:0] out_5813;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5813 (
            .a(out_5812),
            .b(out_3),
            .outp(out_5813)
        );        
        

        logic [WIDTH-1:0] out_5814;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5814 (
            .a(out_5811),
            .b(out_5813),
            .outp(out_5814)
        );        
        

        logic [WIDTH-1:0] out_5815;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5815 (
            .a(out_5808),
            .b(out_5814),
            .outp(out_5815)
        );        
        

        logic [WIDTH-1:0] out_5816;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.05)
        ) inst_5816 (
            .outp(out_5816)
        );
        

        logic [WIDTH-1:0] out_5817;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5817 (
            .a(out_194),
            .b(out_5816),
            .outp(out_5817)
        );        
        

        logic [WIDTH-1:0] out_5818;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5818 (
            .a(out_5442),
            .b(out_5817),
            .outp(out_5818)
        );        
        

        logic [WIDTH-1:0] out_5819;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5)
        ) inst_5819 (
            .outp(out_5819)
        );
        

        logic [WIDTH-1:0] out_5820;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5820 (
            .a(out_5819),
            .b(out_194),
            .outp(out_5820)
        );        
        

        logic [WIDTH-1:0] out_5821;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5821 (
            .a(out_5818),
            .b(out_5820),
            .outp(out_5821)
        );        
        

        logic [WIDTH-1:0] out_5822;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5822 (
            .a(out_14),
            .b(out_4550),
            .outp(out_5822)
        );        
        

        logic [WIDTH-1:0] out_5823;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5823 (
            .in(out_5822),
            .outp(out_5823)
        );
        

        logic [WIDTH-1:0] out_5824;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.3125)
        ) inst_5824 (
            .outp(out_5824)
        );
        

        logic [WIDTH-1:0] out_5825;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5825 (
            .a(out_204),
            .b(out_5824),
            .outp(out_5825)
        );        
        

        logic [WIDTH-1:0] out_5826;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5826 (
            .in(out_5825),
            .outp(out_5826)
        );
        

        logic [WIDTH-1:0] out_5827;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5827 (
            .a(out_5823),
            .b(out_5826),
            .outp(out_5827)
        );        
        

        logic [WIDTH-1:0] out_5828;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5828 (
            .in(out_5827),
            .outp(out_5828)
        );
        

        logic [WIDTH-1:0] out_5829;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5829 (
            .a(out_200),
            .b(out_5828),
            .outp(out_5829)
        );        
        

        logic [WIDTH-1:0] out_5830;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5830 (
            .a(out_5821),
            .b(out_5829),
            .outp(out_5830)
        );        
        

        logic [WIDTH-1:0] out_5831;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5831 (
            .in(out_5817),
            .outp(out_5831)
        );
        

        logic [WIDTH-1:0] out_5832;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5832 (
            .a(out_5823),
            .b(out_5831),
            .outp(out_5832)
        );        
        

        logic [WIDTH-1:0] out_5833;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5833 (
            .in(out_5832),
            .outp(out_5833)
        );
        

        logic [WIDTH-1:0] out_5834;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5834 (
            .a(out_5833),
            .b(out_214),
            .outp(out_5834)
        );        
        

        logic [WIDTH-1:0] out_5835;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5835 (
            .a(out_5830),
            .b(out_5834),
            .outp(out_5835)
        );        
        

        logic [WIDTH-1:0] out_5836;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5836 (
            .a(out_5815),
            .b(out_5835),
            .outp(out_5836)
        );        
        

        logic [WIDTH-1:0] out_5837;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.55)
        ) inst_5837 (
            .outp(out_5837)
        );
        

        logic [WIDTH-1:0] out_5838;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5838 (
            .a(out_5837),
            .b(out_3),
            .outp(out_5838)
        );        
        

        logic [WIDTH-1:0] out_5839;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5839 (
            .in(out_5838),
            .outp(out_5839)
        );
        

        logic [WIDTH-1:0] out_5840;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5840 (
            .a(out_4559),
            .b(out_5839),
            .outp(out_5840)
        );        
        

        logic [WIDTH-1:0] out_5841;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.375)
        ) inst_5841 (
            .outp(out_5841)
        );
        

        logic [WIDTH-1:0] out_5842;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5842 (
            .a(out_5841),
            .b(out_3),
            .outp(out_5842)
        );        
        

        logic [WIDTH-1:0] out_5843;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5843 (
            .a(out_5840),
            .b(out_5842),
            .outp(out_5843)
        );        
        

        logic [WIDTH-1:0] out_5844;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.85)
        ) inst_5844 (
            .outp(out_5844)
        );
        

        logic [WIDTH-1:0] out_5845;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5845 (
            .a(out_5844),
            .b(out_14),
            .outp(out_5845)
        );        
        

        logic [WIDTH-1:0] out_5846;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5846 (
            .a(out_5843),
            .b(out_5845),
            .outp(out_5846)
        );        
        

        logic [WIDTH-1:0] out_5847;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5847 (
            .a(out_5836),
            .b(out_5846),
            .outp(out_5847)
        );        
        

        logic [WIDTH-1:0] out_5848;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5848 (
            .a(out_4551),
            .b(out_5839),
            .outp(out_5848)
        );        
        

        logic [WIDTH-1:0] out_5849;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5)
        ) inst_5849 (
            .outp(out_5849)
        );
        

        logic [WIDTH-1:0] out_5850;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5850 (
            .a(out_14),
            .b(out_5849),
            .outp(out_5850)
        );        
        

        logic [WIDTH-1:0] out_5851;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5851 (
            .a(out_5848),
            .b(out_5850),
            .outp(out_5851)
        );        
        

        logic [WIDTH-1:0] out_5852;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5852 (
            .a(out_5851),
            .b(out_5842),
            .outp(out_5852)
        );        
        

        logic [WIDTH-1:0] out_5853;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5853 (
            .a(out_5847),
            .b(out_5852),
            .outp(out_5853)
        );        
        

        logic [WIDTH-1:0] out_5854;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5854 (
            .a(out_4551),
            .b(out_5800),
            .outp(out_5854)
        );        
        

        logic [WIDTH-1:0] out_5855;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5855 (
            .a(out_5854),
            .b(out_5838),
            .outp(out_5855)
        );        
        

        logic [WIDTH-1:0] out_5856;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.275)
        ) inst_5856 (
            .outp(out_5856)
        );
        

        logic [WIDTH-1:0] out_5857;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5857 (
            .a(out_5856),
            .b(out_3),
            .outp(out_5857)
        );        
        

        logic [WIDTH-1:0] out_5858;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5858 (
            .in(out_5857),
            .outp(out_5858)
        );
        

        logic [WIDTH-1:0] out_5859;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5859 (
            .a(out_5855),
            .b(out_5858),
            .outp(out_5859)
        );        
        

        logic [WIDTH-1:0] out_5860;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5860 (
            .in(out_5839),
            .outp(out_5860)
        );
        

        logic [WIDTH-1:0] out_5861;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5861 (
            .a(out_4534),
            .b(out_5860),
            .outp(out_5861)
        );        
        

        logic [WIDTH-1:0] out_5862;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5862 (
            .in(out_5861),
            .outp(out_5862)
        );
        

        logic [WIDTH-1:0] out_5863;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5863 (
            .a(out_9),
            .b(out_5862),
            .outp(out_5863)
        );        
        

        logic [WIDTH-1:0] out_5864;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5864 (
            .a(out_5859),
            .b(out_5863),
            .outp(out_5864)
        );        
        

        logic [WIDTH-1:0] out_5865;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5865 (
            .a(out_5862),
            .b(out_21),
            .outp(out_5865)
        );        
        

        logic [WIDTH-1:0] out_5866;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5866 (
            .a(out_5864),
            .b(out_5865),
            .outp(out_5866)
        );        
        

        logic [WIDTH-1:0] out_5867;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5867 (
            .a(out_5853),
            .b(out_5866),
            .outp(out_5867)
        );        
        

        logic [WIDTH-1:0] out_5868;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5868 (
            .a(out_1373),
            .b(out_14),
            .outp(out_5868)
        );        
        

        logic [WIDTH-1:0] out_5869;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5869 (
            .a(out_5800),
            .b(out_5868),
            .outp(out_5869)
        );        
        

        logic [WIDTH-1:0] out_5870;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6)
        ) inst_5870 (
            .outp(out_5870)
        );
        

        logic [WIDTH-1:0] out_5871;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5871 (
            .a(out_5870),
            .b(out_3),
            .outp(out_5871)
        );        
        

        logic [WIDTH-1:0] out_5872;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5872 (
            .a(out_5869),
            .b(out_5871),
            .outp(out_5872)
        );        
        

        logic [WIDTH-1:0] out_5873;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5873 (
            .a(out_715),
            .b(out_3),
            .outp(out_5873)
        );        
        

        logic [WIDTH-1:0] out_5874;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5874 (
            .in(out_5873),
            .outp(out_5874)
        );
        

        logic [WIDTH-1:0] out_5875;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5875 (
            .a(out_5872),
            .b(out_5874),
            .outp(out_5875)
        );        
        

        logic [WIDTH-1:0] out_5876;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5876 (
            .a(out_5867),
            .b(out_5875),
            .outp(out_5876)
        );        
        

        logic [WIDTH-1:0] out_5877;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5877 (
            .a(out_4551),
            .b(out_5850),
            .outp(out_5877)
        );        
        

        logic [WIDTH-1:0] out_5878;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5878 (
            .a(out_5877),
            .b(out_5871),
            .outp(out_5878)
        );        
        

        logic [WIDTH-1:0] out_5879;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5879 (
            .a(out_5878),
            .b(out_5874),
            .outp(out_5879)
        );        
        

        logic [WIDTH-1:0] out_5880;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5880 (
            .a(out_5876),
            .b(out_5879),
            .outp(out_5880)
        );        
        

        logic [WIDTH-1:0] out_5881;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5881 (
            .a(out_5434),
            .b(out_4551),
            .outp(out_5881)
        );        
        

        logic [WIDTH-1:0] out_5882;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5882 (
            .a(out_5881),
            .b(out_5800),
            .outp(out_5882)
        );        
        

        logic [WIDTH-1:0] out_5883;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.9)
        ) inst_5883 (
            .outp(out_5883)
        );
        

        logic [WIDTH-1:0] out_5884;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5884 (
            .a(out_5883),
            .b(out_3),
            .outp(out_5884)
        );        
        

        logic [WIDTH-1:0] out_5885;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5885 (
            .in(out_5884),
            .outp(out_5885)
        );
        

        logic [WIDTH-1:0] out_5886;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5886 (
            .a(out_5882),
            .b(out_5885),
            .outp(out_5886)
        );        
        

        logic [WIDTH-1:0] out_5887;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5887 (
            .a(out_5880),
            .b(out_5886),
            .outp(out_5887)
        );        
        

        logic [WIDTH-1:0] out_5888;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1825)
        ) inst_5888 (
            .outp(out_5888)
        );
        

        logic [WIDTH-1:0] out_5889;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5889 (
            .a(out_5888),
            .b(out_127),
            .outp(out_5889)
        );        
        

        logic [WIDTH-1:0] out_5890;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5890 (
            .a(out_5889),
            .b(out_131),
            .outp(out_5890)
        );        
        

        logic [WIDTH-1:0] out_5891;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5891 (
            .a(out_4508),
            .b(out_5890),
            .outp(out_5891)
        );        
        

        logic [WIDTH-1:0] out_5892;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.3775)
        ) inst_5892 (
            .outp(out_5892)
        );
        

        logic [WIDTH-1:0] out_5893;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5893 (
            .a(out_5892),
            .b(out_127),
            .outp(out_5893)
        );        
        

        logic [WIDTH-1:0] out_5894;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5894 (
            .a(out_124),
            .b(out_5893),
            .outp(out_5894)
        );        
        

        logic [WIDTH-1:0] out_5895;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5895 (
            .a(out_5891),
            .b(out_5894),
            .outp(out_5895)
        );        
        

        logic [WIDTH-1:0] out_5896;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5896 (
            .a(out_5887),
            .b(out_5895),
            .outp(out_5896)
        );        
        

        logic [WIDTH-1:0] out_5897;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5897 (
            .a(out_5893),
            .b(out_124),
            .outp(out_5897)
        );        
        

        logic [WIDTH-1:0] out_5898;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5898 (
            .a(out_4513),
            .b(out_5897),
            .outp(out_5898)
        );        
        

        logic [WIDTH-1:0] out_5899;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5899 (
            .a(out_131),
            .b(out_5889),
            .outp(out_5899)
        );        
        

        logic [WIDTH-1:0] out_5900;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5900 (
            .a(out_5898),
            .b(out_5899),
            .outp(out_5900)
        );        
        

        logic [WIDTH-1:0] out_5901;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5901 (
            .a(out_5896),
            .b(out_5900),
            .outp(out_5901)
        );        
        

        logic [WIDTH-1:0] out_5902;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5902 (
            .a(out_4521),
            .b(out_5897),
            .outp(out_5902)
        );        
        

        logic [WIDTH-1:0] out_5903;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.2375)
        ) inst_5903 (
            .outp(out_5903)
        );
        

        logic [WIDTH-1:0] out_5904;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5904 (
            .a(out_5903),
            .b(out_127),
            .outp(out_5904)
        );        
        

        logic [WIDTH-1:0] out_5905;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5905 (
            .a(out_131),
            .b(out_5904),
            .outp(out_5905)
        );        
        

        logic [WIDTH-1:0] out_5906;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5906 (
            .a(out_5902),
            .b(out_5905),
            .outp(out_5906)
        );        
        

        logic [WIDTH-1:0] out_5907;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5907 (
            .a(out_5901),
            .b(out_5906),
            .outp(out_5907)
        );        
        

        logic [WIDTH-1:0] out_5908;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5908 (
            .a(out_4526),
            .b(out_5894),
            .outp(out_5908)
        );        
        

        logic [WIDTH-1:0] out_5909;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5909 (
            .a(out_5904),
            .b(out_131),
            .outp(out_5909)
        );        
        

        logic [WIDTH-1:0] out_5910;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5910 (
            .a(out_5908),
            .b(out_5909),
            .outp(out_5910)
        );        
        

        logic [WIDTH-1:0] out_5911;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5911 (
            .a(out_5907),
            .b(out_5910),
            .outp(out_5911)
        );        
        

        logic [WIDTH-1:0] out_5912;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5375)
        ) inst_5912 (
            .outp(out_5912)
        );
        

        logic [WIDTH-1:0] out_5913;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5913 (
            .a(out_131),
            .b(out_5912),
            .outp(out_5913)
        );        
        

        logic [WIDTH-1:0] out_5914;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5914 (
            .a(out_5913),
            .b(out_127),
            .outp(out_5914)
        );        
        

        logic [WIDTH-1:0] out_5915;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5915 (
            .in(out_5914),
            .outp(out_5915)
        );
        

        logic [WIDTH-1:0] out_5916;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5916 (
            .a(out_4508),
            .b(out_5915),
            .outp(out_5916)
        );        
        

        logic [WIDTH-1:0] out_5917;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.3425)
        ) inst_5917 (
            .outp(out_5917)
        );
        

        logic [WIDTH-1:0] out_5918;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5918 (
            .a(out_5917),
            .b(out_124),
            .outp(out_5918)
        );        
        

        logic [WIDTH-1:0] out_5919;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5919 (
            .a(out_5918),
            .b(out_127),
            .outp(out_5919)
        );        
        

        logic [WIDTH-1:0] out_5920;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5920 (
            .a(out_5916),
            .b(out_5919),
            .outp(out_5920)
        );        
        

        logic [WIDTH-1:0] out_5921;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5921 (
            .a(out_5911),
            .b(out_5920),
            .outp(out_5921)
        );        
        

        logic [WIDTH-1:0] out_5922;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5922 (
            .a(out_4513),
            .b(out_5914),
            .outp(out_5922)
        );        
        

        logic [WIDTH-1:0] out_5923;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5923 (
            .in(out_5919),
            .outp(out_5923)
        );
        

        logic [WIDTH-1:0] out_5924;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5924 (
            .a(out_5922),
            .b(out_5923),
            .outp(out_5924)
        );        
        

        logic [WIDTH-1:0] out_5925;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5925 (
            .a(out_5921),
            .b(out_5924),
            .outp(out_5925)
        );        
        

        logic [WIDTH-1:0] out_5926;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5926 (
            .a(out_4521),
            .b(out_5923),
            .outp(out_5926)
        );        
        

        logic [WIDTH-1:0] out_5927;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.4825)
        ) inst_5927 (
            .outp(out_5927)
        );
        

        logic [WIDTH-1:0] out_5928;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5928 (
            .a(out_131),
            .b(out_5927),
            .outp(out_5928)
        );        
        

        logic [WIDTH-1:0] out_5929;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5929 (
            .a(out_5928),
            .b(out_127),
            .outp(out_5929)
        );        
        

        logic [WIDTH-1:0] out_5930;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5930 (
            .a(out_5926),
            .b(out_5929),
            .outp(out_5930)
        );        
        

        logic [WIDTH-1:0] out_5931;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5931 (
            .a(out_5925),
            .b(out_5930),
            .outp(out_5931)
        );        
        

        logic [WIDTH-1:0] out_5932;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5932 (
            .a(out_4526),
            .b(out_5919),
            .outp(out_5932)
        );        
        

        logic [WIDTH-1:0] out_5933;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5933 (
            .in(out_5929),
            .outp(out_5933)
        );
        

        logic [WIDTH-1:0] out_5934;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5934 (
            .a(out_5932),
            .b(out_5933),
            .outp(out_5934)
        );        
        

        logic [WIDTH-1:0] out_5935;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5935 (
            .a(out_5931),
            .b(out_5934),
            .outp(out_5935)
        );        
        

        logic [WIDTH-1:0] out_5936;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.4575)
        ) inst_5936 (
            .outp(out_5936)
        );
        

        logic [WIDTH-1:0] out_5937;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5937 (
            .a(out_5936),
            .b(out_127),
            .outp(out_5937)
        );        
        

        logic [WIDTH-1:0] out_5938;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5938 (
            .a(out_5937),
            .b(out_131),
            .outp(out_5938)
        );        
        

        logic [WIDTH-1:0] out_5939;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5939 (
            .a(out_4508),
            .b(out_5938),
            .outp(out_5939)
        );        
        

        logic [WIDTH-1:0] out_5940;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6525)
        ) inst_5940 (
            .outp(out_5940)
        );
        

        logic [WIDTH-1:0] out_5941;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5941 (
            .a(out_5940),
            .b(out_127),
            .outp(out_5941)
        );        
        

        logic [WIDTH-1:0] out_5942;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5942 (
            .a(out_124),
            .b(out_5941),
            .outp(out_5942)
        );        
        

        logic [WIDTH-1:0] out_5943;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5943 (
            .a(out_5939),
            .b(out_5942),
            .outp(out_5943)
        );        
        

        logic [WIDTH-1:0] out_5944;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5944 (
            .a(out_5935),
            .b(out_5943),
            .outp(out_5944)
        );        
        

        logic [WIDTH-1:0] out_5945;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5945 (
            .a(out_5941),
            .b(out_124),
            .outp(out_5945)
        );        
        

        logic [WIDTH-1:0] out_5946;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5946 (
            .a(out_4513),
            .b(out_5945),
            .outp(out_5946)
        );        
        

        logic [WIDTH-1:0] out_5947;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5947 (
            .a(out_131),
            .b(out_5937),
            .outp(out_5947)
        );        
        

        logic [WIDTH-1:0] out_5948;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5948 (
            .a(out_5946),
            .b(out_5947),
            .outp(out_5948)
        );        
        

        logic [WIDTH-1:0] out_5949;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5949 (
            .a(out_5944),
            .b(out_5948),
            .outp(out_5949)
        );        
        

        logic [WIDTH-1:0] out_5950;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5950 (
            .a(out_4521),
            .b(out_5945),
            .outp(out_5950)
        );        
        

        logic [WIDTH-1:0] out_5951;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.5125)
        ) inst_5951 (
            .outp(out_5951)
        );
        

        logic [WIDTH-1:0] out_5952;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5952 (
            .a(out_5951),
            .b(out_127),
            .outp(out_5952)
        );        
        

        logic [WIDTH-1:0] out_5953;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5953 (
            .a(out_131),
            .b(out_5952),
            .outp(out_5953)
        );        
        

        logic [WIDTH-1:0] out_5954;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5954 (
            .a(out_5950),
            .b(out_5953),
            .outp(out_5954)
        );        
        

        logic [WIDTH-1:0] out_5955;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5955 (
            .a(out_5949),
            .b(out_5954),
            .outp(out_5955)
        );        
        

        logic [WIDTH-1:0] out_5956;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5956 (
            .a(out_4526),
            .b(out_5942),
            .outp(out_5956)
        );        
        

        logic [WIDTH-1:0] out_5957;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5957 (
            .a(out_5952),
            .b(out_131),
            .outp(out_5957)
        );        
        

        logic [WIDTH-1:0] out_5958;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5958 (
            .a(out_5956),
            .b(out_5957),
            .outp(out_5958)
        );        
        

        logic [WIDTH-1:0] out_5959;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5959 (
            .a(out_5955),
            .b(out_5958),
            .outp(out_5959)
        );        
        

        logic [WIDTH-1:0] out_5960;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.65)
        ) inst_5960 (
            .outp(out_5960)
        );
        

        logic [WIDTH-1:0] out_5961;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5961 (
            .a(out_5960),
            .b(out_14),
            .outp(out_5961)
        );        
        

        logic [WIDTH-1:0] out_5962;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.300001)
        ) inst_5962 (
            .outp(out_5962)
        );
        

        logic [WIDTH-1:0] out_5963;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5963 (
            .a(out_5962),
            .b(out_3),
            .outp(out_5963)
        );        
        

        logic [WIDTH-1:0] out_5964;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5964 (
            .a(out_5961),
            .b(out_5963),
            .outp(out_5964)
        );        
        

        logic [WIDTH-1:0] out_5965;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5965 (
            .a(out_5964),
            .b(out_5800),
            .outp(out_5965)
        );        
        

        logic [WIDTH-1:0] out_5966;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.400001)
        ) inst_5966 (
            .outp(out_5966)
        );
        

        logic [WIDTH-1:0] out_5967;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5967 (
            .a(out_5966),
            .b(out_3),
            .outp(out_5967)
        );        
        

        logic [WIDTH-1:0] out_5968;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5968 (
            .in(out_5967),
            .outp(out_5968)
        );
        

        logic [WIDTH-1:0] out_5969;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5969 (
            .a(out_5965),
            .b(out_5968),
            .outp(out_5969)
        );        
        

        logic [WIDTH-1:0] out_5970;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5970 (
            .a(out_5959),
            .b(out_5969),
            .outp(out_5970)
        );        
        

        logic [WIDTH-1:0] out_5971;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5971 (
            .a(out_3505),
            .b(out_5510),
            .outp(out_5971)
        );        
        

        logic [WIDTH-1:0] out_5972;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5972 (
            .a(out_4558),
            .b(out_14),
            .outp(out_5972)
        );        
        

        logic [WIDTH-1:0] out_5973;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5973 (
            .a(out_5971),
            .b(out_5972),
            .outp(out_5973)
        );        
        

        logic [WIDTH-1:0] out_5974;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.550001)
        ) inst_5974 (
            .outp(out_5974)
        );
        

        logic [WIDTH-1:0] out_5975;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5975 (
            .a(out_5974),
            .b(out_3),
            .outp(out_5975)
        );        
        

        logic [WIDTH-1:0] out_5976;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5976 (
            .in(out_5975),
            .outp(out_5976)
        );
        

        logic [WIDTH-1:0] out_5977;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5977 (
            .a(out_5973),
            .b(out_5976),
            .outp(out_5977)
        );        
        

        logic [WIDTH-1:0] out_5978;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5978 (
            .a(out_5970),
            .b(out_5977),
            .outp(out_5978)
        );        
        

        logic [WIDTH-1:0] out_5979;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5979 (
            .a(out_3505),
            .b(out_4551),
            .outp(out_5979)
        );        
        

        logic [WIDTH-1:0] out_5980;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5980 (
            .a(out_5979),
            .b(out_5976),
            .outp(out_5980)
        );        
        

        logic [WIDTH-1:0] out_5981;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5981 (
            .a(out_14),
            .b(out_5960),
            .outp(out_5981)
        );        
        

        logic [WIDTH-1:0] out_5982;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5982 (
            .a(out_5980),
            .b(out_5981),
            .outp(out_5982)
        );        
        

        logic [WIDTH-1:0] out_5983;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5983 (
            .in(out_5981),
            .outp(out_5983)
        );
        

        logic [WIDTH-1:0] out_5984;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5984 (
            .a(out_3506),
            .b(out_5983),
            .outp(out_5984)
        );        
        

        logic [WIDTH-1:0] out_5985;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5985 (
            .in(out_5984),
            .outp(out_5985)
        );
        

        logic [WIDTH-1:0] out_5986;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5986 (
            .a(out_336),
            .b(out_5985),
            .outp(out_5986)
        );        
        

        logic [WIDTH-1:0] out_5987;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5987 (
            .a(out_5982),
            .b(out_5986),
            .outp(out_5987)
        );        
        

        logic [WIDTH-1:0] out_5988;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5988 (
            .a(out_5985),
            .b(out_343),
            .outp(out_5988)
        );        
        

        logic [WIDTH-1:0] out_5989;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5989 (
            .a(out_5987),
            .b(out_5988),
            .outp(out_5989)
        );        
        

        logic [WIDTH-1:0] out_5990;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5990 (
            .a(out_5978),
            .b(out_5989),
            .outp(out_5990)
        );        
        

        logic [WIDTH-1:0] out_5991;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.65875)
        ) inst_5991 (
            .outp(out_5991)
        );
        

        logic [WIDTH-1:0] out_5992;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5992 (
            .a(out_5991),
            .b(out_1891),
            .outp(out_5992)
        );        
        

        logic [WIDTH-1:0] out_5993;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5993 (
            .a(out_5992),
            .b(out_137),
            .outp(out_5993)
        );        
        

        logic [WIDTH-1:0] out_5994;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.281875)
        ) inst_5994 (
            .outp(out_5994)
        );
        

        logic [WIDTH-1:0] out_5995;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5995 (
            .a(out_5994),
            .b(out_4052),
            .outp(out_5995)
        );        
        

        logic [WIDTH-1:0] out_5996;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5996 (
            .a(out_5993),
            .b(out_5995),
            .outp(out_5996)
        );        
        

        logic [WIDTH-1:0] out_5997;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.13813)
        ) inst_5997 (
            .outp(out_5997)
        );
        

        logic [WIDTH-1:0] out_5998;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5998 (
            .a(out_1907),
            .b(out_5997),
            .outp(out_5998)
        );        
        

        logic [WIDTH-1:0] out_5999;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_5999 (
            .a(out_1904),
            .b(out_5998),
            .outp(out_5999)
        );        
        

        logic [WIDTH-1:0] out_6000;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6000 (
            .a(out_5996),
            .b(out_5999),
            .outp(out_6000)
        );        
        

        logic [WIDTH-1:0] out_6001;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.13813)
        ) inst_6001 (
            .outp(out_6001)
        );
        

        logic [WIDTH-1:0] out_6002;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6002 (
            .a(out_1907),
            .b(out_6001),
            .outp(out_6002)
        );        
        

        logic [WIDTH-1:0] out_6003;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6003 (
            .a(out_6002),
            .b(out_1904),
            .outp(out_6003)
        );        
        

        logic [WIDTH-1:0] out_6004;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6004 (
            .a(out_4052),
            .b(out_5994),
            .outp(out_6004)
        );        
        

        logic [WIDTH-1:0] out_6005;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6005 (
            .a(out_6003),
            .b(out_6004),
            .outp(out_6005)
        );        
        

        logic [WIDTH-1:0] out_6006;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6006 (
            .a(out_137),
            .b(out_5992),
            .outp(out_6006)
        );        
        

        logic [WIDTH-1:0] out_6007;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6007 (
            .a(out_6005),
            .b(out_6006),
            .outp(out_6007)
        );        
        

        logic [WIDTH-1:0] out_6008;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6008 (
            .a(out_6000),
            .b(out_6007),
            .outp(out_6008)
        );        
        

        logic [WIDTH-1:0] out_6009;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6009 (
            .in(out_6008),
            .outp(out_6009)
        );
        

        logic [WIDTH-1:0] out_6010;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.475)
        ) inst_6010 (
            .outp(out_6010)
        );
        

        logic [WIDTH-1:0] out_6011;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6011 (
            .a(out_14),
            .b(out_6010),
            .outp(out_6011)
        );        
        

        logic [WIDTH-1:0] out_6012;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6012 (
            .a(out_6009),
            .b(out_6011),
            .outp(out_6012)
        );        
        

        logic [WIDTH-1:0] out_6013;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.25)
        ) inst_6013 (
            .outp(out_6013)
        );
        

        logic [WIDTH-1:0] out_6014;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6014 (
            .a(out_6013),
            .b(out_14),
            .outp(out_6014)
        );        
        

        logic [WIDTH-1:0] out_6015;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6015 (
            .a(out_6012),
            .b(out_6014),
            .outp(out_6015)
        );        
        

        logic [WIDTH-1:0] out_6016;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.375)
        ) inst_6016 (
            .outp(out_6016)
        );
        

        logic [WIDTH-1:0] out_6017;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6017 (
            .a(out_6016),
            .b(out_3),
            .outp(out_6017)
        );        
        

        logic [WIDTH-1:0] out_6018;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6018 (
            .a(out_6015),
            .b(out_6017),
            .outp(out_6018)
        );        
        

        logic [WIDTH-1:0] out_6019;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.525)
        ) inst_6019 (
            .outp(out_6019)
        );
        

        logic [WIDTH-1:0] out_6020;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6020 (
            .a(out_6019),
            .b(out_3),
            .outp(out_6020)
        );        
        

        logic [WIDTH-1:0] out_6021;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6021 (
            .in(out_6020),
            .outp(out_6021)
        );
        

        logic [WIDTH-1:0] out_6022;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6022 (
            .a(out_6018),
            .b(out_6021),
            .outp(out_6022)
        );        
        

        logic [WIDTH-1:0] out_6023;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.491667)
        ) inst_6023 (
            .outp(out_6023)
        );
        

        logic [WIDTH-1:0] out_6024;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6024 (
            .a(out_1933),
            .b(out_6023),
            .outp(out_6024)
        );        
        

        logic [WIDTH-1:0] out_6025;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6025 (
            .in(out_6024),
            .outp(out_6025)
        );
        

        logic [WIDTH-1:0] out_6026;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.45)
        ) inst_6026 (
            .outp(out_6026)
        );
        

        logic [WIDTH-1:0] out_6027;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6027 (
            .a(out_6026),
            .b(out_3),
            .outp(out_6027)
        );        
        

        logic [WIDTH-1:0] out_6028;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6028 (
            .in(out_6027),
            .outp(out_6028)
        );
        

        logic [WIDTH-1:0] out_6029;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6029 (
            .a(out_6025),
            .b(out_6028),
            .outp(out_6029)
        );        
        

        logic [WIDTH-1:0] out_6030;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6030 (
            .in(out_6029),
            .outp(out_6030)
        );
        

        logic [WIDTH-1:0] out_6031;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6031 (
            .a(out_6030),
            .b(out_460),
            .outp(out_6031)
        );        
        

        logic [WIDTH-1:0] out_6032;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6032 (
            .a(out_6022),
            .b(out_6031),
            .outp(out_6032)
        );        
        

        logic [WIDTH-1:0] out_6033;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6033 (
            .a(out_5990),
            .b(out_6032),
            .outp(out_6033)
        );        
        

        logic [WIDTH-1:0] out_6034;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6034 (
            .in(out_6011),
            .outp(out_6034)
        );
        

        logic [WIDTH-1:0] out_6035;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.425)
        ) inst_6035 (
            .outp(out_6035)
        );
        

        logic [WIDTH-1:0] out_6036;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6036 (
            .a(out_6035),
            .b(out_3),
            .outp(out_6036)
        );        
        

        logic [WIDTH-1:0] out_6037;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6037 (
            .in(out_6036),
            .outp(out_6037)
        );
        

        logic [WIDTH-1:0] out_6038;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6038 (
            .a(out_6034),
            .b(out_6037),
            .outp(out_6038)
        );        
        

        logic [WIDTH-1:0] out_6039;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6039 (
            .in(out_6038),
            .outp(out_6039)
        );
        

        logic [WIDTH-1:0] out_6040;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6040 (
            .a(out_6039),
            .b(out_460),
            .outp(out_6040)
        );        
        

        logic [WIDTH-1:0] out_6041;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6041 (
            .a(out_6033),
            .b(out_6040),
            .outp(out_6041)
        );        
        

        logic [WIDTH-1:0] out_6042;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.9)
        ) inst_6042 (
            .outp(out_6042)
        );
        

        logic [WIDTH-1:0] out_6043;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6043 (
            .a(out_6042),
            .b(out_3),
            .outp(out_6043)
        );        
        

        logic [WIDTH-1:0] out_6044;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6044 (
            .in(out_6043),
            .outp(out_6044)
        );
        

        logic [WIDTH-1:0] out_6045;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6045 (
            .a(out_4534),
            .b(out_6044),
            .outp(out_6045)
        );        
        

        logic [WIDTH-1:0] out_6046;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6046 (
            .in(out_6045),
            .outp(out_6046)
        );
        

        logic [WIDTH-1:0] out_6047;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6047 (
            .a(out_9),
            .b(out_6046),
            .outp(out_6047)
        );        
        

        logic [WIDTH-1:0] out_6048;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6048 (
            .a(out_6046),
            .b(out_21),
            .outp(out_6048)
        );        
        

        logic [WIDTH-1:0] out_6049;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6049 (
            .a(out_6047),
            .b(out_6048),
            .outp(out_6049)
        );        
        

        logic [WIDTH-1:0] out_6050;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6050 (
            .a(out_6041),
            .b(out_6049),
            .outp(out_6050)
        );        
        

        logic [WIDTH-1:0] out_6051;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6051 (
            .in(out_5842),
            .outp(out_6051)
        );
        

        logic [WIDTH-1:0] out_6052;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6052 (
            .a(out_5854),
            .b(out_6051),
            .outp(out_6052)
        );        
        

        logic [WIDTH-1:0] out_6053;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.275)
        ) inst_6053 (
            .outp(out_6053)
        );
        

        logic [WIDTH-1:0] out_6054;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6054 (
            .a(out_6053),
            .b(out_3),
            .outp(out_6054)
        );        
        

        logic [WIDTH-1:0] out_6055;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6055 (
            .a(out_6052),
            .b(out_6054),
            .outp(out_6055)
        );        
        

        logic [WIDTH-1:0] out_6056;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6056 (
            .a(out_6050),
            .b(out_6055),
            .outp(out_6056)
        );        
        

        logic [WIDTH-1:0] out_6057;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.951)
        ) inst_6057 (
            .outp(out_6057)
        );
        

        logic [WIDTH-1:0] out_6058;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6058 (
            .a(out_3),
            .b(out_6057),
            .outp(out_6058)
        );        
        

        logic [WIDTH-1:0] out_6059;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6059 (
            .in(out_6058),
            .outp(out_6059)
        );
        

        logic [WIDTH-1:0] out_6060;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6060 (
            .a(out_14),
            .b(out_252),
            .outp(out_6060)
        );        
        

        logic [WIDTH-1:0] out_6061;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6061 (
            .in(out_6060),
            .outp(out_6061)
        );
        

        logic [WIDTH-1:0] out_6062;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6062 (
            .a(out_6059),
            .b(out_6061),
            .outp(out_6062)
        );        
        

        logic [WIDTH-1:0] out_6063;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6063 (
            .in(out_6062),
            .outp(out_6063)
        );
        

        logic [WIDTH-1:0] out_6064;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6064 (
            .a(out_6063),
            .b(out_21),
            .outp(out_6064)
        );        
        

        logic [WIDTH-1:0] out_6065;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.226)
        ) inst_6065 (
            .outp(out_6065)
        );
        

        logic [WIDTH-1:0] out_6066;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6066 (
            .a(out_3),
            .b(out_6065),
            .outp(out_6066)
        );        
        

        logic [WIDTH-1:0] out_6067;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6067 (
            .a(out_6064),
            .b(out_6066),
            .outp(out_6067)
        );        
        

        logic [WIDTH-1:0] out_6068;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.676)
        ) inst_6068 (
            .outp(out_6068)
        );
        

        logic [WIDTH-1:0] out_6069;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6069 (
            .a(out_6068),
            .b(out_3),
            .outp(out_6069)
        );        
        

        logic [WIDTH-1:0] out_6070;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6070 (
            .a(out_6067),
            .b(out_6069),
            .outp(out_6070)
        );        
        

        logic [WIDTH-1:0] out_6071;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6071 (
            .a(out_9),
            .b(out_6063),
            .outp(out_6071)
        );        
        

        logic [WIDTH-1:0] out_6072;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6072 (
            .a(out_6070),
            .b(out_6071),
            .outp(out_6072)
        );        
        

        logic [WIDTH-1:0] out_6073;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.25)
        ) inst_6073 (
            .outp(out_6073)
        );
        

        logic [WIDTH-1:0] out_6074;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6074 (
            .a(out_14),
            .b(out_6073),
            .outp(out_6074)
        );        
        

        logic [WIDTH-1:0] out_6075;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6075 (
            .a(out_6072),
            .b(out_6074),
            .outp(out_6075)
        );        
        

        logic [WIDTH-1:0] out_6076;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.025)
        ) inst_6076 (
            .outp(out_6076)
        );
        

        logic [WIDTH-1:0] out_6077;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6077 (
            .a(out_6076),
            .b(out_14),
            .outp(out_6077)
        );        
        

        logic [WIDTH-1:0] out_6078;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6078 (
            .a(out_6075),
            .b(out_6077),
            .outp(out_6078)
        );        
        

        logic [WIDTH-1:0] out_6079;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6079 (
            .a(out_6056),
            .b(out_6078),
            .outp(out_6079)
        );        
        

        logic [WIDTH-1:0] out_6080;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.05)
        ) inst_6080 (
            .outp(out_6080)
        );
        

        logic [WIDTH-1:0] out_6081;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6081 (
            .a(out_14),
            .b(out_6080),
            .outp(out_6081)
        );        
        

        logic [WIDTH-1:0] out_6082;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.556)
        ) inst_6082 (
            .outp(out_6082)
        );
        

        logic [WIDTH-1:0] out_6083;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6083 (
            .a(out_3),
            .b(out_6082),
            .outp(out_6083)
        );        
        

        logic [WIDTH-1:0] out_6084;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6084 (
            .a(out_6081),
            .b(out_6083),
            .outp(out_6084)
        );        
        

        logic [WIDTH-1:0] out_6085;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.456)
        ) inst_6085 (
            .outp(out_6085)
        );
        

        logic [WIDTH-1:0] out_6086;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6086 (
            .a(out_6085),
            .b(out_3),
            .outp(out_6086)
        );        
        

        logic [WIDTH-1:0] out_6087;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6087 (
            .a(out_6084),
            .b(out_6086),
            .outp(out_6087)
        );        
        

        logic [WIDTH-1:0] out_6088;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6088 (
            .a(out_66),
            .b(out_14),
            .outp(out_6088)
        );        
        

        logic [WIDTH-1:0] out_6089;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6089 (
            .a(out_6087),
            .b(out_6088),
            .outp(out_6089)
        );        
        

        logic [WIDTH-1:0] out_6090;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6090 (
            .a(out_6079),
            .b(out_6089),
            .outp(out_6090)
        );        
        

        logic [WIDTH-1:0] out_6091;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.146856)
        ) inst_6091 (
            .outp(out_6091)
        );
        

        logic [WIDTH-1:0] out_6092;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6092 (
            .a(out_6091),
            .b(out_3),
            .outp(out_6092)
        );        
        

        logic [WIDTH-1:0] out_6093;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6093 (
            .a(out_6092),
            .b(out_1495),
            .outp(out_6093)
        );        
        

        logic [WIDTH-1:0] out_6094;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6094 (
            .in(out_6093),
            .outp(out_6094)
        );
        

        logic [WIDTH-1:0] out_6095;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6095 (
            .a(out_6094),
            .b(out_6061),
            .outp(out_6095)
        );        
        

        logic [WIDTH-1:0] out_6096;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6096 (
            .in(out_6095),
            .outp(out_6096)
        );
        

        logic [WIDTH-1:0] out_6097;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6097 (
            .a(out_9),
            .b(out_6096),
            .outp(out_6097)
        );        
        

        logic [WIDTH-1:0] out_6098;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6098 (
            .a(out_6096),
            .b(out_21),
            .outp(out_6098)
        );        
        

        logic [WIDTH-1:0] out_6099;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6099 (
            .a(out_6097),
            .b(out_6098),
            .outp(out_6099)
        );        
        

        logic [WIDTH-1:0] out_6100;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6100 (
            .a(out_6090),
            .b(out_6099),
            .outp(out_6100)
        );        
        

        logic [WIDTH-1:0] out_6101;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.44765)
        ) inst_6101 (
            .outp(out_6101)
        );
        

        logic [WIDTH-1:0] out_6102;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6102 (
            .a(out_6101),
            .b(out_1891),
            .outp(out_6102)
        );        
        

        logic [WIDTH-1:0] out_6103;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6103 (
            .a(out_6102),
            .b(out_137),
            .outp(out_6103)
        );        
        

        logic [WIDTH-1:0] out_6104;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.27973)
        ) inst_6104 (
            .outp(out_6104)
        );
        

        logic [WIDTH-1:0] out_6105;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6105 (
            .a(out_6104),
            .b(out_4052),
            .outp(out_6105)
        );        
        

        logic [WIDTH-1:0] out_6106;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6106 (
            .a(out_6103),
            .b(out_6105),
            .outp(out_6106)
        );        
        

        logic [WIDTH-1:0] out_6107;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.92488)
        ) inst_6107 (
            .outp(out_6107)
        );
        

        logic [WIDTH-1:0] out_6108;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6108 (
            .a(out_1907),
            .b(out_6107),
            .outp(out_6108)
        );        
        

        logic [WIDTH-1:0] out_6109;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6109 (
            .a(out_1904),
            .b(out_6108),
            .outp(out_6109)
        );        
        

        logic [WIDTH-1:0] out_6110;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6110 (
            .a(out_6106),
            .b(out_6109),
            .outp(out_6110)
        );        
        

        logic [WIDTH-1:0] out_6111;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6111 (
            .a(out_6108),
            .b(out_1904),
            .outp(out_6111)
        );        
        

        logic [WIDTH-1:0] out_6112;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6112 (
            .a(out_4052),
            .b(out_6104),
            .outp(out_6112)
        );        
        

        logic [WIDTH-1:0] out_6113;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6113 (
            .a(out_6111),
            .b(out_6112),
            .outp(out_6113)
        );        
        

        logic [WIDTH-1:0] out_6114;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6114 (
            .a(out_137),
            .b(out_6102),
            .outp(out_6114)
        );        
        

        logic [WIDTH-1:0] out_6115;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6115 (
            .a(out_6113),
            .b(out_6114),
            .outp(out_6115)
        );        
        

        logic [WIDTH-1:0] out_6116;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6116 (
            .a(out_6110),
            .b(out_6115),
            .outp(out_6116)
        );        
        

        logic [WIDTH-1:0] out_6117;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6117 (
            .in(out_6116),
            .outp(out_6117)
        );
        

        logic [WIDTH-1:0] out_6118;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.775)
        ) inst_6118 (
            .outp(out_6118)
        );
        

        logic [WIDTH-1:0] out_6119;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6119 (
            .a(out_14),
            .b(out_6118),
            .outp(out_6119)
        );        
        

        logic [WIDTH-1:0] out_6120;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6120 (
            .a(out_6117),
            .b(out_6119),
            .outp(out_6120)
        );        
        

        logic [WIDTH-1:0] out_6121;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.55)
        ) inst_6121 (
            .outp(out_6121)
        );
        

        logic [WIDTH-1:0] out_6122;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6122 (
            .a(out_6121),
            .b(out_14),
            .outp(out_6122)
        );        
        

        logic [WIDTH-1:0] out_6123;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6123 (
            .a(out_6120),
            .b(out_6122),
            .outp(out_6123)
        );        
        

        logic [WIDTH-1:0] out_6124;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.171)
        ) inst_6124 (
            .outp(out_6124)
        );
        

        logic [WIDTH-1:0] out_6125;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6125 (
            .a(out_3),
            .b(out_6124),
            .outp(out_6125)
        );        
        

        logic [WIDTH-1:0] out_6126;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6126 (
            .a(out_6123),
            .b(out_6125),
            .outp(out_6126)
        );        
        

        logic [WIDTH-1:0] out_6127;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0209999)
        ) inst_6127 (
            .outp(out_6127)
        );
        

        logic [WIDTH-1:0] out_6128;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6128 (
            .a(out_6127),
            .b(out_3),
            .outp(out_6128)
        );        
        

        logic [WIDTH-1:0] out_6129;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6129 (
            .a(out_6126),
            .b(out_6128),
            .outp(out_6129)
        );        
        

        logic [WIDTH-1:0] out_6130;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.59167)
        ) inst_6130 (
            .outp(out_6130)
        );
        

        logic [WIDTH-1:0] out_6131;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6131 (
            .a(out_1933),
            .b(out_6130),
            .outp(out_6131)
        );        
        

        logic [WIDTH-1:0] out_6132;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6132 (
            .in(out_6131),
            .outp(out_6132)
        );
        

        logic [WIDTH-1:0] out_6133;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0959997)
        ) inst_6133 (
            .outp(out_6133)
        );
        

        logic [WIDTH-1:0] out_6134;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6134 (
            .a(out_3),
            .b(out_6133),
            .outp(out_6134)
        );        
        

        logic [WIDTH-1:0] out_6135;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6135 (
            .in(out_6134),
            .outp(out_6135)
        );
        

        logic [WIDTH-1:0] out_6136;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6136 (
            .a(out_6132),
            .b(out_6135),
            .outp(out_6136)
        );        
        

        logic [WIDTH-1:0] out_6137;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6137 (
            .in(out_6136),
            .outp(out_6137)
        );
        

        logic [WIDTH-1:0] out_6138;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6138 (
            .a(out_6137),
            .b(out_460),
            .outp(out_6138)
        );        
        

        logic [WIDTH-1:0] out_6139;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6139 (
            .a(out_6129),
            .b(out_6138),
            .outp(out_6139)
        );        
        

        logic [WIDTH-1:0] out_6140;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6140 (
            .a(out_6100),
            .b(out_6139),
            .outp(out_6140)
        );        
        

        logic [WIDTH-1:0] out_6141;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6141 (
            .in(out_6119),
            .outp(out_6141)
        );
        

        logic [WIDTH-1:0] out_6142;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.121)
        ) inst_6142 (
            .outp(out_6142)
        );
        

        logic [WIDTH-1:0] out_6143;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6143 (
            .a(out_3),
            .b(out_6142),
            .outp(out_6143)
        );        
        

        logic [WIDTH-1:0] out_6144;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6144 (
            .in(out_6143),
            .outp(out_6144)
        );
        

        logic [WIDTH-1:0] out_6145;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6145 (
            .a(out_6141),
            .b(out_6144),
            .outp(out_6145)
        );        
        

        logic [WIDTH-1:0] out_6146;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6146 (
            .in(out_6145),
            .outp(out_6146)
        );
        

        logic [WIDTH-1:0] out_6147;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6147 (
            .a(out_6146),
            .b(out_460),
            .outp(out_6147)
        );        
        

        logic [WIDTH-1:0] out_6148;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6148 (
            .a(out_6140),
            .b(out_6147),
            .outp(out_6148)
        );        
        

        logic [WIDTH-1:0] out_6149;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.525)
        ) inst_6149 (
            .outp(out_6149)
        );
        

        logic [WIDTH-1:0] out_6150;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6150 (
            .a(out_6149),
            .b(out_137),
            .outp(out_6150)
        );        
        

        logic [WIDTH-1:0] out_6151;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.12055)
        ) inst_6151 (
            .outp(out_6151)
        );
        

        logic [WIDTH-1:0] out_6152;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6152 (
            .a(out_4480),
            .b(out_6151),
            .outp(out_6152)
        );        
        

        logic [WIDTH-1:0] out_6153;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6153 (
            .a(out_6150),
            .b(out_6152),
            .outp(out_6153)
        );        
        

        logic [WIDTH-1:0] out_6154;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.65055)
        ) inst_6154 (
            .outp(out_6154)
        );
        

        logic [WIDTH-1:0] out_6155;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6155 (
            .a(out_6154),
            .b(out_4477),
            .outp(out_6155)
        );        
        

        logic [WIDTH-1:0] out_6156;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6156 (
            .a(out_6153),
            .b(out_6155),
            .outp(out_6156)
        );        
        

        logic [WIDTH-1:0] out_6157;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6157 (
            .a(out_6148),
            .b(out_6156),
            .outp(out_6157)
        );        
        

        logic [WIDTH-1:0] out_6158;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.02555)
        ) inst_6158 (
            .outp(out_6158)
        );
        

        logic [WIDTH-1:0] out_6159;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6159 (
            .a(out_6158),
            .b(out_131),
            .outp(out_6159)
        );        
        

        logic [WIDTH-1:0] out_6160;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6160 (
            .a(out_127),
            .b(out_6159),
            .outp(out_6160)
        );        
        

        logic [WIDTH-1:0] out_6161;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.500551)
        ) inst_6161 (
            .outp(out_6161)
        );
        

        logic [WIDTH-1:0] out_6162;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6162 (
            .a(out_6161),
            .b(out_124),
            .outp(out_6162)
        );        
        

        logic [WIDTH-1:0] out_6163;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6163 (
            .a(out_6162),
            .b(out_127),
            .outp(out_6163)
        );        
        

        logic [WIDTH-1:0] out_6164;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6164 (
            .a(out_6160),
            .b(out_6163),
            .outp(out_6164)
        );        
        

        logic [WIDTH-1:0] out_6165;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.47)
        ) inst_6165 (
            .outp(out_6165)
        );
        

        logic [WIDTH-1:0] out_6166;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6166 (
            .a(out_6165),
            .b(out_152),
            .outp(out_6166)
        );        
        

        logic [WIDTH-1:0] out_6167;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6167 (
            .a(out_6164),
            .b(out_6166),
            .outp(out_6167)
        );        
        

        logic [WIDTH-1:0] out_6168;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6168 (
            .a(out_6157),
            .b(out_6167),
            .outp(out_6168)
        );        
        

        logic [WIDTH-1:0] out_6169;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6169 (
            .a(out_127),
            .b(out_6162),
            .outp(out_6169)
        );        
        

        logic [WIDTH-1:0] out_6170;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6170 (
            .a(out_6159),
            .b(out_127),
            .outp(out_6170)
        );        
        

        logic [WIDTH-1:0] out_6171;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6171 (
            .a(out_6169),
            .b(out_6170),
            .outp(out_6171)
        );        
        

        logic [WIDTH-1:0] out_6172;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6172 (
            .a(out_152),
            .b(out_6165),
            .outp(out_6172)
        );        
        

        logic [WIDTH-1:0] out_6173;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6173 (
            .a(out_6171),
            .b(out_6172),
            .outp(out_6173)
        );        
        

        logic [WIDTH-1:0] out_6174;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6174 (
            .a(out_6168),
            .b(out_6173),
            .outp(out_6174)
        );        
        

        logic [WIDTH-1:0] out_6175;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.970551)
        ) inst_6175 (
            .outp(out_6175)
        );
        

        logic [WIDTH-1:0] out_6176;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6176 (
            .a(out_6175),
            .b(out_131),
            .outp(out_6176)
        );        
        

        logic [WIDTH-1:0] out_6177;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6177 (
            .a(out_6176),
            .b(out_127),
            .outp(out_6177)
        );        
        

        logic [WIDTH-1:0] out_6178;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6178 (
            .a(out_6169),
            .b(out_6177),
            .outp(out_6178)
        );        
        

        logic [WIDTH-1:0] out_6179;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6179 (
            .a(out_137),
            .b(out_6149),
            .outp(out_6179)
        );        
        

        logic [WIDTH-1:0] out_6180;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6180 (
            .a(out_6178),
            .b(out_6179),
            .outp(out_6180)
        );        
        

        logic [WIDTH-1:0] out_6181;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6181 (
            .a(out_6174),
            .b(out_6180),
            .outp(out_6181)
        );        
        

        logic [WIDTH-1:0] out_6182;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.970552)
        ) inst_6182 (
            .outp(out_6182)
        );
        

        logic [WIDTH-1:0] out_6183;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6183 (
            .a(out_6182),
            .b(out_131),
            .outp(out_6183)
        );        
        

        logic [WIDTH-1:0] out_6184;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6184 (
            .a(out_127),
            .b(out_6183),
            .outp(out_6184)
        );        
        

        logic [WIDTH-1:0] out_6185;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6185 (
            .a(out_6163),
            .b(out_6184),
            .outp(out_6185)
        );        
        

        logic [WIDTH-1:0] out_6186;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6186 (
            .a(out_6185),
            .b(out_6150),
            .outp(out_6186)
        );        
        

        logic [WIDTH-1:0] out_6187;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6187 (
            .a(out_6181),
            .b(out_6186),
            .outp(out_6187)
        );        
        

        logic [WIDTH-1:0] out_6188;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.32055)
        ) inst_6188 (
            .outp(out_6188)
        );
        

        logic [WIDTH-1:0] out_6189;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6189 (
            .a(out_6188),
            .b(out_4477),
            .outp(out_6189)
        );        
        

        logic [WIDTH-1:0] out_6190;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.84555)
        ) inst_6190 (
            .outp(out_6190)
        );
        

        logic [WIDTH-1:0] out_6191;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6191 (
            .a(out_4480),
            .b(out_6190),
            .outp(out_6191)
        );        
        

        logic [WIDTH-1:0] out_6192;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6192 (
            .a(out_6189),
            .b(out_6191),
            .outp(out_6192)
        );        
        

        logic [WIDTH-1:0] out_6193;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6193 (
            .a(out_6192),
            .b(out_6166),
            .outp(out_6193)
        );        
        

        logic [WIDTH-1:0] out_6194;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6194 (
            .a(out_6187),
            .b(out_6193),
            .outp(out_6194)
        );        
        

        logic [WIDTH-1:0] out_6195;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6195 (
            .a(out_6190),
            .b(out_4480),
            .outp(out_6195)
        );        
        

        logic [WIDTH-1:0] out_6196;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6196 (
            .a(out_4477),
            .b(out_6188),
            .outp(out_6196)
        );        
        

        logic [WIDTH-1:0] out_6197;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6197 (
            .a(out_6195),
            .b(out_6196),
            .outp(out_6197)
        );        
        

        logic [WIDTH-1:0] out_6198;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6198 (
            .a(out_6197),
            .b(out_6172),
            .outp(out_6198)
        );        
        

        logic [WIDTH-1:0] out_6199;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6199 (
            .a(out_6194),
            .b(out_6198),
            .outp(out_6199)
        );        
        

        logic [WIDTH-1:0] out_6200;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.37555)
        ) inst_6200 (
            .outp(out_6200)
        );
        

        logic [WIDTH-1:0] out_6201;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6201 (
            .a(out_4477),
            .b(out_6200),
            .outp(out_6201)
        );        
        

        logic [WIDTH-1:0] out_6202;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6202 (
            .a(out_6195),
            .b(out_6201),
            .outp(out_6202)
        );        
        

        logic [WIDTH-1:0] out_6203;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6203 (
            .a(out_6202),
            .b(out_6179),
            .outp(out_6203)
        );        
        

        logic [WIDTH-1:0] out_6204;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6204 (
            .a(out_6199),
            .b(out_6203),
            .outp(out_6204)
        );        
        

        logic [WIDTH-1:0] out_6205;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.37555)
        ) inst_6205 (
            .outp(out_6205)
        );
        

        logic [WIDTH-1:0] out_6206;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6206 (
            .a(out_6205),
            .b(out_4477),
            .outp(out_6206)
        );        
        

        logic [WIDTH-1:0] out_6207;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6207 (
            .a(out_6191),
            .b(out_6206),
            .outp(out_6207)
        );        
        

        logic [WIDTH-1:0] out_6208;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6208 (
            .a(out_6207),
            .b(out_6150),
            .outp(out_6208)
        );        
        

        logic [WIDTH-1:0] out_6209;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6209 (
            .a(out_6204),
            .b(out_6208),
            .outp(out_6209)
        );        
        

        logic [WIDTH-1:0] out_6210;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.751)
        ) inst_6210 (
            .outp(out_6210)
        );
        

        logic [WIDTH-1:0] out_6211;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6211 (
            .a(out_6210),
            .b(out_3),
            .outp(out_6211)
        );        
        

        logic [WIDTH-1:0] out_6212;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.851)
        ) inst_6212 (
            .outp(out_6212)
        );
        

        logic [WIDTH-1:0] out_6213;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6213 (
            .a(out_3),
            .b(out_6212),
            .outp(out_6213)
        );        
        

        logic [WIDTH-1:0] out_6214;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6214 (
            .a(out_6211),
            .b(out_6213),
            .outp(out_6214)
        );        
        

        logic [WIDTH-1:0] out_6215;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.7)
        ) inst_6215 (
            .outp(out_6215)
        );
        

        logic [WIDTH-1:0] out_6216;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6216 (
            .a(out_14),
            .b(out_6215),
            .outp(out_6216)
        );        
        

        logic [WIDTH-1:0] out_6217;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6217 (
            .a(out_6214),
            .b(out_6216),
            .outp(out_6217)
        );        
        

        logic [WIDTH-1:0] out_6218;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6218 (
            .a(out_6217),
            .b(out_6088),
            .outp(out_6218)
        );        
        

        logic [WIDTH-1:0] out_6219;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6219 (
            .a(out_6209),
            .b(out_6218),
            .outp(out_6219)
        );        
        

        logic [WIDTH-1:0] out_6220;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6220 (
            .a(out_680),
            .b(out_14),
            .outp(out_6220)
        );        
        

        logic [WIDTH-1:0] out_6221;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.576)
        ) inst_6221 (
            .outp(out_6221)
        );
        

        logic [WIDTH-1:0] out_6222;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6222 (
            .a(out_6221),
            .b(out_3),
            .outp(out_6222)
        );        
        

        logic [WIDTH-1:0] out_6223;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6223 (
            .a(out_6220),
            .b(out_6222),
            .outp(out_6223)
        );        
        

        logic [WIDTH-1:0] out_6224;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.751)
        ) inst_6224 (
            .outp(out_6224)
        );
        

        logic [WIDTH-1:0] out_6225;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6225 (
            .a(out_3),
            .b(out_6224),
            .outp(out_6225)
        );        
        

        logic [WIDTH-1:0] out_6226;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6226 (
            .a(out_6223),
            .b(out_6225),
            .outp(out_6226)
        );        
        

        logic [WIDTH-1:0] out_6227;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6227 (
            .a(out_6226),
            .b(out_6074),
            .outp(out_6227)
        );        
        

        logic [WIDTH-1:0] out_6228;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6228 (
            .a(out_6219),
            .b(out_6227),
            .outp(out_6228)
        );        
        

        logic [WIDTH-1:0] out_6229;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6229 (
            .a(out_6222),
            .b(out_6225),
            .outp(out_6229)
        );        
        

        logic [WIDTH-1:0] out_6230;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.8)
        ) inst_6230 (
            .outp(out_6230)
        );
        

        logic [WIDTH-1:0] out_6231;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6231 (
            .a(out_14),
            .b(out_6230),
            .outp(out_6231)
        );        
        

        logic [WIDTH-1:0] out_6232;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6232 (
            .a(out_6229),
            .b(out_6231),
            .outp(out_6232)
        );        
        

        logic [WIDTH-1:0] out_6233;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6233 (
            .a(out_6232),
            .b(out_6088),
            .outp(out_6233)
        );        
        

        logic [WIDTH-1:0] out_6234;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6234 (
            .a(out_6228),
            .b(out_6233),
            .outp(out_6234)
        );        
        

        logic [WIDTH-1:0] out_6235;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.851)
        ) inst_6235 (
            .outp(out_6235)
        );
        

        logic [WIDTH-1:0] out_6236;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6236 (
            .a(out_6235),
            .b(out_3),
            .outp(out_6236)
        );        
        

        logic [WIDTH-1:0] out_6237;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.576)
        ) inst_6237 (
            .outp(out_6237)
        );
        

        logic [WIDTH-1:0] out_6238;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6238 (
            .a(out_3),
            .b(out_6237),
            .outp(out_6238)
        );        
        

        logic [WIDTH-1:0] out_6239;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6239 (
            .a(out_6236),
            .b(out_6238),
            .outp(out_6239)
        );        
        

        logic [WIDTH-1:0] out_6240;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6240 (
            .in(out_6222),
            .outp(out_6240)
        );
        

        logic [WIDTH-1:0] out_6241;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6241 (
            .a(out_6240),
            .b(out_6061),
            .outp(out_6241)
        );        
        

        logic [WIDTH-1:0] out_6242;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6242 (
            .in(out_6241),
            .outp(out_6242)
        );
        

        logic [WIDTH-1:0] out_6243;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6243 (
            .a(out_9),
            .b(out_6242),
            .outp(out_6243)
        );        
        

        logic [WIDTH-1:0] out_6244;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6244 (
            .a(out_6239),
            .b(out_6243),
            .outp(out_6244)
        );        
        

        logic [WIDTH-1:0] out_6245;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6245 (
            .a(out_6242),
            .b(out_21),
            .outp(out_6245)
        );        
        

        logic [WIDTH-1:0] out_6246;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6246 (
            .a(out_6244),
            .b(out_6245),
            .outp(out_6246)
        );        
        

        logic [WIDTH-1:0] out_6247;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6247 (
            .a(out_6246),
            .b(out_6216),
            .outp(out_6247)
        );        
        

        logic [WIDTH-1:0] out_6248;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6248 (
            .a(out_6247),
            .b(out_6088),
            .outp(out_6248)
        );        
        

        logic [WIDTH-1:0] out_6249;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6249 (
            .a(out_6234),
            .b(out_6248),
            .outp(out_6249)
        );        
        

        logic [WIDTH-1:0] out_6250;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.126)
        ) inst_6250 (
            .outp(out_6250)
        );
        

        logic [WIDTH-1:0] out_6251;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6251 (
            .a(out_6250),
            .b(out_3),
            .outp(out_6251)
        );        
        

        logic [WIDTH-1:0] out_6252;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6252 (
            .a(out_6066),
            .b(out_6251),
            .outp(out_6252)
        );        
        

        logic [WIDTH-1:0] out_6253;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6253 (
            .a(out_14),
            .b(out_6076),
            .outp(out_6253)
        );        
        

        logic [WIDTH-1:0] out_6254;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6254 (
            .a(out_6252),
            .b(out_6253),
            .outp(out_6254)
        );        
        

        logic [WIDTH-1:0] out_6255;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6255 (
            .a(out_6254),
            .b(out_6088),
            .outp(out_6255)
        );        
        

        logic [WIDTH-1:0] out_6256;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6256 (
            .a(out_6249),
            .b(out_6255),
            .outp(out_6256)
        );        
        

        logic [WIDTH-1:0] out_6257;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.776)
        ) inst_6257 (
            .outp(out_6257)
        );
        

        logic [WIDTH-1:0] out_6258;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6258 (
            .a(out_3),
            .b(out_6257),
            .outp(out_6258)
        );        
        

        logic [WIDTH-1:0] out_6259;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6259 (
            .a(out_6258),
            .b(out_6069),
            .outp(out_6259)
        );        
        

        logic [WIDTH-1:0] out_6260;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6260 (
            .a(out_6259),
            .b(out_6088),
            .outp(out_6260)
        );        
        

        logic [WIDTH-1:0] out_6261;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6261 (
            .a(out_6260),
            .b(out_6074),
            .outp(out_6261)
        );        
        

        logic [WIDTH-1:0] out_6262;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6262 (
            .a(out_6256),
            .b(out_6261),
            .outp(out_6262)
        );        
        

        logic [WIDTH-1:0] out_6263;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6263 (
            .a(out_58),
            .b(out_14),
            .outp(out_6263)
        );        
        

        logic [WIDTH-1:0] out_6264;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.862)
        ) inst_6264 (
            .outp(out_6264)
        );
        

        logic [WIDTH-1:0] out_6265;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6265 (
            .a(out_6264),
            .b(out_3),
            .outp(out_6265)
        );        
        

        logic [WIDTH-1:0] out_6266;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6266 (
            .a(out_6263),
            .b(out_6265),
            .outp(out_6266)
        );        
        

        logic [WIDTH-1:0] out_6267;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.962)
        ) inst_6267 (
            .outp(out_6267)
        );
        

        logic [WIDTH-1:0] out_6268;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6268 (
            .a(out_6267),
            .b(out_3),
            .outp(out_6268)
        );        
        

        logic [WIDTH-1:0] out_6269;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6269 (
            .in(out_6268),
            .outp(out_6269)
        );
        

        logic [WIDTH-1:0] out_6270;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6270 (
            .a(out_6266),
            .b(out_6269),
            .outp(out_6270)
        );        
        

        logic [WIDTH-1:0] out_6271;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6271 (
            .a(out_6270),
            .b(out_6074),
            .outp(out_6271)
        );        
        

        logic [WIDTH-1:0] out_6272;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6272 (
            .a(out_6262),
            .b(out_6271),
            .outp(out_6272)
        );        
        

        logic [WIDTH-1:0] out_6273;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.4)
        ) inst_6273 (
            .outp(out_6273)
        );
        

        logic [WIDTH-1:0] out_6274;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6274 (
            .a(out_14),
            .b(out_6273),
            .outp(out_6274)
        );        
        

        logic [WIDTH-1:0] out_6275;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6275 (
            .in(out_6274),
            .outp(out_6275)
        );
        

        logic [WIDTH-1:0] out_6276;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.912)
        ) inst_6276 (
            .outp(out_6276)
        );
        

        logic [WIDTH-1:0] out_6277;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6277 (
            .a(out_6276),
            .b(out_3),
            .outp(out_6277)
        );        
        

        logic [WIDTH-1:0] out_6278;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6278 (
            .in(out_6277),
            .outp(out_6278)
        );
        

        logic [WIDTH-1:0] out_6279;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6279 (
            .a(out_6275),
            .b(out_6278),
            .outp(out_6279)
        );        
        

        logic [WIDTH-1:0] out_6280;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6280 (
            .in(out_6279),
            .outp(out_6280)
        );
        

        logic [WIDTH-1:0] out_6281;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6281 (
            .a(out_6280),
            .b(out_460),
            .outp(out_6281)
        );        
        

        logic [WIDTH-1:0] out_6282;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6282 (
            .a(out_6272),
            .b(out_6281),
            .outp(out_6282)
        );        
        

        logic [WIDTH-1:0] out_6283;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.662)
        ) inst_6283 (
            .outp(out_6283)
        );
        

        logic [WIDTH-1:0] out_6284;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6284 (
            .a(out_6283),
            .b(out_3),
            .outp(out_6284)
        );        
        

        logic [WIDTH-1:0] out_6285;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.762)
        ) inst_6285 (
            .outp(out_6285)
        );
        

        logic [WIDTH-1:0] out_6286;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6286 (
            .a(out_6285),
            .b(out_3),
            .outp(out_6286)
        );        
        

        logic [WIDTH-1:0] out_6287;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6287 (
            .in(out_6286),
            .outp(out_6287)
        );
        

        logic [WIDTH-1:0] out_6288;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6288 (
            .a(out_6284),
            .b(out_6287),
            .outp(out_6288)
        );        
        

        logic [WIDTH-1:0] out_6289;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6289 (
            .a(out_6288),
            .b(out_6216),
            .outp(out_6289)
        );        
        

        logic [WIDTH-1:0] out_6290;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6290 (
            .a(out_6289),
            .b(out_6088),
            .outp(out_6290)
        );        
        

        logic [WIDTH-1:0] out_6291;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6291 (
            .a(out_6282),
            .b(out_6290),
            .outp(out_6291)
        );        
        

        logic [WIDTH-1:0] out_6292;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.487)
        ) inst_6292 (
            .outp(out_6292)
        );
        

        logic [WIDTH-1:0] out_6293;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6293 (
            .a(out_6292),
            .b(out_3),
            .outp(out_6293)
        );        
        

        logic [WIDTH-1:0] out_6294;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6294 (
            .a(out_6220),
            .b(out_6293),
            .outp(out_6294)
        );        
        

        logic [WIDTH-1:0] out_6295;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6295 (
            .in(out_6284),
            .outp(out_6295)
        );
        

        logic [WIDTH-1:0] out_6296;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6296 (
            .a(out_6294),
            .b(out_6295),
            .outp(out_6296)
        );        
        

        logic [WIDTH-1:0] out_6297;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6297 (
            .a(out_6296),
            .b(out_6074),
            .outp(out_6297)
        );        
        

        logic [WIDTH-1:0] out_6298;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6298 (
            .a(out_6291),
            .b(out_6297),
            .outp(out_6298)
        );        
        

        logic [WIDTH-1:0] out_6299;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6299 (
            .a(out_6231),
            .b(out_6293),
            .outp(out_6299)
        );        
        

        logic [WIDTH-1:0] out_6300;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6300 (
            .a(out_6299),
            .b(out_6295),
            .outp(out_6300)
        );        
        

        logic [WIDTH-1:0] out_6301;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6301 (
            .a(out_6300),
            .b(out_6088),
            .outp(out_6301)
        );        
        

        logic [WIDTH-1:0] out_6302;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6302 (
            .a(out_6298),
            .b(out_6301),
            .outp(out_6302)
        );        
        

        logic [WIDTH-1:0] out_6303;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.762)
        ) inst_6303 (
            .outp(out_6303)
        );
        

        logic [WIDTH-1:0] out_6304;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6304 (
            .a(out_6303),
            .b(out_3),
            .outp(out_6304)
        );        
        

        logic [WIDTH-1:0] out_6305;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6305 (
            .in(out_6293),
            .outp(out_6305)
        );
        

        logic [WIDTH-1:0] out_6306;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6306 (
            .a(out_6304),
            .b(out_6305),
            .outp(out_6306)
        );        
        

        logic [WIDTH-1:0] out_6307;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6307 (
            .in(out_6293),
            .outp(out_6307)
        );
        

        logic [WIDTH-1:0] out_6308;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6308 (
            .a(out_6307),
            .b(out_6061),
            .outp(out_6308)
        );        
        

        logic [WIDTH-1:0] out_6309;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6309 (
            .in(out_6308),
            .outp(out_6309)
        );
        

        logic [WIDTH-1:0] out_6310;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6310 (
            .a(out_9),
            .b(out_6309),
            .outp(out_6310)
        );        
        

        logic [WIDTH-1:0] out_6311;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6311 (
            .a(out_6306),
            .b(out_6310),
            .outp(out_6311)
        );        
        

        logic [WIDTH-1:0] out_6312;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6312 (
            .a(out_6309),
            .b(out_21),
            .outp(out_6312)
        );        
        

        logic [WIDTH-1:0] out_6313;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6313 (
            .a(out_6311),
            .b(out_6312),
            .outp(out_6313)
        );        
        

        logic [WIDTH-1:0] out_6314;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6314 (
            .a(out_6313),
            .b(out_6216),
            .outp(out_6314)
        );        
        

        logic [WIDTH-1:0] out_6315;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6315 (
            .a(out_6314),
            .b(out_6088),
            .outp(out_6315)
        );        
        

        logic [WIDTH-1:0] out_6316;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6316 (
            .a(out_6302),
            .b(out_6315),
            .outp(out_6316)
        );        
        

        logic [WIDTH-1:0] out_6317;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.882)
        ) inst_6317 (
            .outp(out_6317)
        );
        

        logic [WIDTH-1:0] out_6318;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6318 (
            .a(out_6317),
            .b(out_3),
            .outp(out_6318)
        );        
        

        logic [WIDTH-1:0] out_6319;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6319 (
            .a(out_6081),
            .b(out_6318),
            .outp(out_6319)
        );        
        

        logic [WIDTH-1:0] out_6320;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.982)
        ) inst_6320 (
            .outp(out_6320)
        );
        

        logic [WIDTH-1:0] out_6321;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6321 (
            .a(out_6320),
            .b(out_3),
            .outp(out_6321)
        );        
        

        logic [WIDTH-1:0] out_6322;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6322 (
            .in(out_6321),
            .outp(out_6322)
        );
        

        logic [WIDTH-1:0] out_6323;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6323 (
            .a(out_6319),
            .b(out_6322),
            .outp(out_6323)
        );        
        

        logic [WIDTH-1:0] out_6324;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6324 (
            .a(out_6323),
            .b(out_6088),
            .outp(out_6324)
        );        
        

        logic [WIDTH-1:0] out_6325;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6325 (
            .a(out_6316),
            .b(out_6324),
            .outp(out_6325)
        );        
        

        logic [WIDTH-1:0] out_6326;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.58486)
        ) inst_6326 (
            .outp(out_6326)
        );
        

        logic [WIDTH-1:0] out_6327;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6327 (
            .a(out_6326),
            .b(out_3),
            .outp(out_6327)
        );        
        

        logic [WIDTH-1:0] out_6328;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6328 (
            .a(out_6327),
            .b(out_1495),
            .outp(out_6328)
        );        
        

        logic [WIDTH-1:0] out_6329;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6329 (
            .in(out_6328),
            .outp(out_6329)
        );
        

        logic [WIDTH-1:0] out_6330;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6330 (
            .a(out_6329),
            .b(out_6061),
            .outp(out_6330)
        );        
        

        logic [WIDTH-1:0] out_6331;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6331 (
            .in(out_6330),
            .outp(out_6331)
        );
        

        logic [WIDTH-1:0] out_6332;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6332 (
            .a(out_9),
            .b(out_6331),
            .outp(out_6332)
        );        
        

        logic [WIDTH-1:0] out_6333;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6333 (
            .a(out_6331),
            .b(out_21),
            .outp(out_6333)
        );        
        

        logic [WIDTH-1:0] out_6334;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6334 (
            .a(out_6332),
            .b(out_6333),
            .outp(out_6334)
        );        
        

        logic [WIDTH-1:0] out_6335;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6335 (
            .a(out_6325),
            .b(out_6334),
            .outp(out_6335)
        );        
        

        logic [WIDTH-1:0] out_6336;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0790005)
        ) inst_6336 (
            .outp(out_6336)
        );
        

        logic [WIDTH-1:0] out_6337;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6337 (
            .a(out_6336),
            .b(out_3),
            .outp(out_6337)
        );        
        

        logic [WIDTH-1:0] out_6338;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.579001)
        ) inst_6338 (
            .outp(out_6338)
        );
        

        logic [WIDTH-1:0] out_6339;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6339 (
            .a(out_6338),
            .b(out_3),
            .outp(out_6339)
        );        
        

        logic [WIDTH-1:0] out_6340;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6340 (
            .in(out_6339),
            .outp(out_6340)
        );
        

        logic [WIDTH-1:0] out_6341;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6341 (
            .a(out_6337),
            .b(out_6340),
            .outp(out_6341)
        );        
        

        logic [WIDTH-1:0] out_6342;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.015)
        ) inst_6342 (
            .outp(out_6342)
        );
        

        logic [WIDTH-1:0] out_6343;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6343 (
            .a(out_14),
            .b(out_6342),
            .outp(out_6343)
        );        
        

        logic [WIDTH-1:0] out_6344;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6344 (
            .a(out_6341),
            .b(out_6343),
            .outp(out_6344)
        );        
        

        logic [WIDTH-1:0] out_6345;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6345 (
            .a(out_684),
            .b(out_14),
            .outp(out_6345)
        );        
        

        logic [WIDTH-1:0] out_6346;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6346 (
            .a(out_6344),
            .b(out_6345),
            .outp(out_6346)
        );        
        

        logic [WIDTH-1:0] out_6347;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.354001)
        ) inst_6347 (
            .outp(out_6347)
        );
        

        logic [WIDTH-1:0] out_6348;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6348 (
            .a(out_6347),
            .b(out_3),
            .outp(out_6348)
        );        
        

        logic [WIDTH-1:0] out_6349;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6349 (
            .in(out_6348),
            .outp(out_6349)
        );
        

        logic [WIDTH-1:0] out_6350;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6350 (
            .a(out_6349),
            .b(out_6061),
            .outp(out_6350)
        );        
        

        logic [WIDTH-1:0] out_6351;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6351 (
            .in(out_6350),
            .outp(out_6351)
        );
        

        logic [WIDTH-1:0] out_6352;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6352 (
            .a(out_6351),
            .b(out_21),
            .outp(out_6352)
        );        
        

        logic [WIDTH-1:0] out_6353;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.712975)
        ) inst_6353 (
            .outp(out_6353)
        );
        

        logic [WIDTH-1:0] out_6354;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6354 (
            .a(out_6353),
            .b(out_556),
            .outp(out_6354)
        );        
        

        logic [WIDTH-1:0] out_6355;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6355 (
            .a(out_6354),
            .b(out_559),
            .outp(out_6355)
        );        
        

        logic [WIDTH-1:0] out_6356;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.34202)
        ) inst_6356 (
            .outp(out_6356)
        );
        

        logic [WIDTH-1:0] out_6357;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6357 (
            .a(out_6356),
            .b(out_2653),
            .outp(out_6357)
        );        
        

        logic [WIDTH-1:0] out_6358;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6358 (
            .a(out_6355),
            .b(out_6357),
            .outp(out_6358)
        );        
        

        logic [WIDTH-1:0] out_6359;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.23375)
        ) inst_6359 (
            .outp(out_6359)
        );
        

        logic [WIDTH-1:0] out_6360;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6360 (
            .a(out_553),
            .b(out_6359),
            .outp(out_6360)
        );        
        

        logic [WIDTH-1:0] out_6361;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6361 (
            .a(out_6358),
            .b(out_6360),
            .outp(out_6361)
        );        
        

        logic [WIDTH-1:0] out_6362;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6362 (
            .a(out_2653),
            .b(out_6356),
            .outp(out_6362)
        );        
        

        logic [WIDTH-1:0] out_6363;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6363 (
            .a(out_559),
            .b(out_6354),
            .outp(out_6363)
        );        
        

        logic [WIDTH-1:0] out_6364;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6364 (
            .a(out_6362),
            .b(out_6363),
            .outp(out_6364)
        );        
        

        logic [WIDTH-1:0] out_6365;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6365 (
            .a(out_6359),
            .b(out_553),
            .outp(out_6365)
        );        
        

        logic [WIDTH-1:0] out_6366;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6366 (
            .a(out_6364),
            .b(out_6365),
            .outp(out_6366)
        );        
        

        logic [WIDTH-1:0] out_6367;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6367 (
            .a(out_6361),
            .b(out_6366),
            .outp(out_6367)
        );        
        

        logic [WIDTH-1:0] out_6368;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6368 (
            .in(out_6367),
            .outp(out_6368)
        );
        

        logic [WIDTH-1:0] out_6369;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6369 (
            .a(out_6352),
            .b(out_6368),
            .outp(out_6369)
        );        
        

        logic [WIDTH-1:0] out_6370;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6370 (
            .a(out_9),
            .b(out_6351),
            .outp(out_6370)
        );        
        

        logic [WIDTH-1:0] out_6371;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6371 (
            .a(out_6369),
            .b(out_6370),
            .outp(out_6371)
        );        
        

        logic [WIDTH-1:0] out_6372;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6372 (
            .a(out_6346),
            .b(out_6371),
            .outp(out_6372)
        );        
        

        logic [WIDTH-1:0] out_6373;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6373 (
            .a(out_6352),
            .b(out_6372),
            .outp(out_6373)
        );        
        

        logic [WIDTH-1:0] out_6374;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6374 (
            .a(out_6335),
            .b(out_6373),
            .outp(out_6374)
        );        
        

        logic [WIDTH-1:0] out_6375;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.987)
        ) inst_6375 (
            .outp(out_6375)
        );
        

        logic [WIDTH-1:0] out_6376;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6376 (
            .a(out_6375),
            .b(out_3),
            .outp(out_6376)
        );        
        

        logic [WIDTH-1:0] out_6377;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.087)
        ) inst_6377 (
            .outp(out_6377)
        );
        

        logic [WIDTH-1:0] out_6378;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6378 (
            .a(out_6377),
            .b(out_3),
            .outp(out_6378)
        );        
        

        logic [WIDTH-1:0] out_6379;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6379 (
            .in(out_6378),
            .outp(out_6379)
        );
        

        logic [WIDTH-1:0] out_6380;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6380 (
            .a(out_6376),
            .b(out_6379),
            .outp(out_6380)
        );        
        

        logic [WIDTH-1:0] out_6381;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6381 (
            .a(out_6380),
            .b(out_6088),
            .outp(out_6381)
        );        
        

        logic [WIDTH-1:0] out_6382;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6382 (
            .a(out_6381),
            .b(out_6074),
            .outp(out_6382)
        );        
        

        logic [WIDTH-1:0] out_6383;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6383 (
            .a(out_6374),
            .b(out_6382),
            .outp(out_6383)
        );        
        

        logic [WIDTH-1:0] out_6384;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.00286)
        ) inst_6384 (
            .outp(out_6384)
        );
        

        logic [WIDTH-1:0] out_6385;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6385 (
            .a(out_6384),
            .b(out_194),
            .outp(out_6385)
        );        
        

        logic [WIDTH-1:0] out_6386;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.55286)
        ) inst_6386 (
            .outp(out_6386)
        );
        

        logic [WIDTH-1:0] out_6387;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6387 (
            .a(out_6386),
            .b(out_194),
            .outp(out_6387)
        );        
        

        logic [WIDTH-1:0] out_6388;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6388 (
            .in(out_6387),
            .outp(out_6388)
        );
        

        logic [WIDTH-1:0] out_6389;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6389 (
            .a(out_6385),
            .b(out_6388),
            .outp(out_6389)
        );        
        

        logic [WIDTH-1:0] out_6390;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6390 (
            .a(out_14),
            .b(out_66),
            .outp(out_6390)
        );        
        

        logic [WIDTH-1:0] out_6391;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6391 (
            .in(out_6390),
            .outp(out_6391)
        );
        

        logic [WIDTH-1:0] out_6392;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.25357)
        ) inst_6392 (
            .outp(out_6392)
        );
        

        logic [WIDTH-1:0] out_6393;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6393 (
            .a(out_6392),
            .b(out_204),
            .outp(out_6393)
        );        
        

        logic [WIDTH-1:0] out_6394;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6394 (
            .in(out_6393),
            .outp(out_6394)
        );
        

        logic [WIDTH-1:0] out_6395;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6395 (
            .a(out_6391),
            .b(out_6394),
            .outp(out_6395)
        );        
        

        logic [WIDTH-1:0] out_6396;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6396 (
            .in(out_6395),
            .outp(out_6396)
        );
        

        logic [WIDTH-1:0] out_6397;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6397 (
            .a(out_200),
            .b(out_6396),
            .outp(out_6397)
        );        
        

        logic [WIDTH-1:0] out_6398;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6398 (
            .a(out_6389),
            .b(out_6397),
            .outp(out_6398)
        );        
        

        logic [WIDTH-1:0] out_6399;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6399 (
            .in(out_6385),
            .outp(out_6399)
        );
        

        logic [WIDTH-1:0] out_6400;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6400 (
            .a(out_6391),
            .b(out_6399),
            .outp(out_6400)
        );        
        

        logic [WIDTH-1:0] out_6401;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6401 (
            .in(out_6400),
            .outp(out_6401)
        );
        

        logic [WIDTH-1:0] out_6402;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6402 (
            .a(out_6401),
            .b(out_214),
            .outp(out_6402)
        );        
        

        logic [WIDTH-1:0] out_6403;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6403 (
            .a(out_6398),
            .b(out_6402),
            .outp(out_6403)
        );        
        

        logic [WIDTH-1:0] out_6404;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6404 (
            .a(out_6403),
            .b(out_6088),
            .outp(out_6404)
        );        
        

        logic [WIDTH-1:0] out_6405;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6405 (
            .a(out_6404),
            .b(out_6074),
            .outp(out_6405)
        );        
        

        logic [WIDTH-1:0] out_6406;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6406 (
            .a(out_6383),
            .b(out_6405),
            .outp(out_6406)
        );        
        

        logic [WIDTH-1:0] out_6407;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.187)
        ) inst_6407 (
            .outp(out_6407)
        );
        

        logic [WIDTH-1:0] out_6408;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6408 (
            .a(out_6407),
            .b(out_3),
            .outp(out_6408)
        );        
        

        logic [WIDTH-1:0] out_6409;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.287)
        ) inst_6409 (
            .outp(out_6409)
        );
        

        logic [WIDTH-1:0] out_6410;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6410 (
            .a(out_6409),
            .b(out_3),
            .outp(out_6410)
        );        
        

        logic [WIDTH-1:0] out_6411;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6411 (
            .in(out_6410),
            .outp(out_6411)
        );
        

        logic [WIDTH-1:0] out_6412;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6412 (
            .a(out_6408),
            .b(out_6411),
            .outp(out_6412)
        );        
        

        logic [WIDTH-1:0] out_6413;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6413 (
            .a(out_6412),
            .b(out_6088),
            .outp(out_6413)
        );        
        

        logic [WIDTH-1:0] out_6414;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6414 (
            .a(out_6413),
            .b(out_6074),
            .outp(out_6414)
        );        
        

        logic [WIDTH-1:0] out_6415;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6415 (
            .a(out_6406),
            .b(out_6414),
            .outp(out_6415)
        );        
        

        logic [WIDTH-1:0] out_6416;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.637)
        ) inst_6416 (
            .outp(out_6416)
        );
        

        logic [WIDTH-1:0] out_6417;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6417 (
            .a(out_6416),
            .b(out_3),
            .outp(out_6417)
        );        
        

        logic [WIDTH-1:0] out_6418;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.737)
        ) inst_6418 (
            .outp(out_6418)
        );
        

        logic [WIDTH-1:0] out_6419;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6419 (
            .a(out_6418),
            .b(out_3),
            .outp(out_6419)
        );        
        

        logic [WIDTH-1:0] out_6420;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6420 (
            .in(out_6419),
            .outp(out_6420)
        );
        

        logic [WIDTH-1:0] out_6421;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6421 (
            .a(out_6417),
            .b(out_6420),
            .outp(out_6421)
        );        
        

        logic [WIDTH-1:0] out_6422;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6422 (
            .a(out_252),
            .b(out_14),
            .outp(out_6422)
        );        
        

        logic [WIDTH-1:0] out_6423;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6423 (
            .a(out_6421),
            .b(out_6422),
            .outp(out_6423)
        );        
        

        logic [WIDTH-1:0] out_6424;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6424 (
            .a(out_6423),
            .b(out_6074),
            .outp(out_6424)
        );        
        

        logic [WIDTH-1:0] out_6425;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6425 (
            .a(out_6415),
            .b(out_6424),
            .outp(out_6425)
        );        
        

        logic [WIDTH-1:0] out_6426;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6426 (
            .a(out_6408),
            .b(out_6420),
            .outp(out_6426)
        );        
        

        logic [WIDTH-1:0] out_6427;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.462)
        ) inst_6427 (
            .outp(out_6427)
        );
        

        logic [WIDTH-1:0] out_6428;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6428 (
            .a(out_6427),
            .b(out_3),
            .outp(out_6428)
        );        
        

        logic [WIDTH-1:0] out_6429;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6429 (
            .in(out_6428),
            .outp(out_6429)
        );
        

        logic [WIDTH-1:0] out_6430;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6430 (
            .a(out_6429),
            .b(out_6061),
            .outp(out_6430)
        );        
        

        logic [WIDTH-1:0] out_6431;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6431 (
            .in(out_6430),
            .outp(out_6431)
        );
        

        logic [WIDTH-1:0] out_6432;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6432 (
            .a(out_9),
            .b(out_6431),
            .outp(out_6432)
        );        
        

        logic [WIDTH-1:0] out_6433;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6433 (
            .a(out_6426),
            .b(out_6432),
            .outp(out_6433)
        );        
        

        logic [WIDTH-1:0] out_6434;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6434 (
            .a(out_6431),
            .b(out_21),
            .outp(out_6434)
        );        
        

        logic [WIDTH-1:0] out_6435;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6435 (
            .a(out_6433),
            .b(out_6434),
            .outp(out_6435)
        );        
        

        logic [WIDTH-1:0] out_6436;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6436 (
            .a(out_6435),
            .b(out_6088),
            .outp(out_6436)
        );        
        

        logic [WIDTH-1:0] out_6437;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6437 (
            .a(out_6436),
            .b(out_6060),
            .outp(out_6437)
        );        
        

        logic [WIDTH-1:0] out_6438;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6438 (
            .a(out_6425),
            .b(out_6437),
            .outp(out_6438)
        );        
        

        logic [WIDTH-1:0] out_6439;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.325)
        ) inst_6439 (
            .outp(out_6439)
        );
        

        logic [WIDTH-1:0] out_6440;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6440 (
            .a(out_6439),
            .b(out_14),
            .outp(out_6440)
        );        
        

        logic [WIDTH-1:0] out_6441;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.587)
        ) inst_6441 (
            .outp(out_6441)
        );
        

        logic [WIDTH-1:0] out_6442;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6442 (
            .a(out_6441),
            .b(out_3),
            .outp(out_6442)
        );        
        

        logic [WIDTH-1:0] out_6443;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6443 (
            .a(out_6440),
            .b(out_6442),
            .outp(out_6443)
        );        
        

        logic [WIDTH-1:0] out_6444;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.137)
        ) inst_6444 (
            .outp(out_6444)
        );
        

        logic [WIDTH-1:0] out_6445;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6445 (
            .a(out_6444),
            .b(out_3),
            .outp(out_6445)
        );        
        

        logic [WIDTH-1:0] out_6446;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6446 (
            .in(out_6445),
            .outp(out_6446)
        );
        

        logic [WIDTH-1:0] out_6447;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6447 (
            .a(out_6443),
            .b(out_6446),
            .outp(out_6447)
        );        
        

        logic [WIDTH-1:0] out_6448;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6448 (
            .a(out_14),
            .b(out_58),
            .outp(out_6448)
        );        
        

        logic [WIDTH-1:0] out_6449;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6449 (
            .in(out_6448),
            .outp(out_6449)
        );
        

        logic [WIDTH-1:0] out_6450;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6450 (
            .in(out_6445),
            .outp(out_6450)
        );
        

        logic [WIDTH-1:0] out_6451;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6451 (
            .a(out_6449),
            .b(out_6450),
            .outp(out_6451)
        );        
        

        logic [WIDTH-1:0] out_6452;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6452 (
            .in(out_6451),
            .outp(out_6452)
        );
        

        logic [WIDTH-1:0] out_6453;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6453 (
            .a(out_9),
            .b(out_6452),
            .outp(out_6453)
        );        
        

        logic [WIDTH-1:0] out_6454;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6454 (
            .a(out_6447),
            .b(out_6453),
            .outp(out_6454)
        );        
        

        logic [WIDTH-1:0] out_6455;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6455 (
            .a(out_6452),
            .b(out_21),
            .outp(out_6455)
        );        
        

        logic [WIDTH-1:0] out_6456;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6456 (
            .a(out_6454),
            .b(out_6455),
            .outp(out_6456)
        );        
        

        logic [WIDTH-1:0] out_6457;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6457 (
            .a(out_6456),
            .b(out_6448),
            .outp(out_6457)
        );        
        

        logic [WIDTH-1:0] out_6458;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6458 (
            .a(out_6438),
            .b(out_6457),
            .outp(out_6458)
        );        
        

        logic [WIDTH-1:0] out_6459;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.9)
        ) inst_6459 (
            .outp(out_6459)
        );
        

        logic [WIDTH-1:0] out_6460;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6460 (
            .a(out_14),
            .b(out_6459),
            .outp(out_6460)
        );        
        

        logic [WIDTH-1:0] out_6461;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.8)
        ) inst_6461 (
            .outp(out_6461)
        );
        

        logic [WIDTH-1:0] out_6462;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6462 (
            .a(out_6461),
            .b(out_14),
            .outp(out_6462)
        );        
        

        logic [WIDTH-1:0] out_6463;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6463 (
            .a(out_6460),
            .b(out_6462),
            .outp(out_6463)
        );        
        

        logic [WIDTH-1:0] out_6464;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.5305)
        ) inst_6464 (
            .outp(out_6464)
        );
        

        logic [WIDTH-1:0] out_6465;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6465 (
            .a(out_3),
            .b(out_6464),
            .outp(out_6465)
        );        
        

        logic [WIDTH-1:0] out_6466;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6466 (
            .a(out_6463),
            .b(out_6465),
            .outp(out_6466)
        );        
        

        logic [WIDTH-1:0] out_6467;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.0305)
        ) inst_6467 (
            .outp(out_6467)
        );
        

        logic [WIDTH-1:0] out_6468;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6468 (
            .a(out_6467),
            .b(out_3),
            .outp(out_6468)
        );        
        

        logic [WIDTH-1:0] out_6469;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6469 (
            .a(out_6466),
            .b(out_6468),
            .outp(out_6469)
        );        
        

        logic [WIDTH-1:0] out_6470;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6470 (
            .a(out_6458),
            .b(out_6469),
            .outp(out_6470)
        );        
        

        logic [WIDTH-1:0] out_6471;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.3305)
        ) inst_6471 (
            .outp(out_6471)
        );
        

        logic [WIDTH-1:0] out_6472;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6472 (
            .a(out_3),
            .b(out_6471),
            .outp(out_6472)
        );        
        

        logic [WIDTH-1:0] out_6473;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6473 (
            .a(out_6462),
            .b(out_6472),
            .outp(out_6473)
        );        
        

        logic [WIDTH-1:0] out_6474;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.2305)
        ) inst_6474 (
            .outp(out_6474)
        );
        

        logic [WIDTH-1:0] out_6475;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6475 (
            .a(out_6474),
            .b(out_3),
            .outp(out_6475)
        );        
        

        logic [WIDTH-1:0] out_6476;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6476 (
            .a(out_6473),
            .b(out_6475),
            .outp(out_6476)
        );        
        

        logic [WIDTH-1:0] out_6477;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6477 (
            .a(out_14),
            .b(out_3043),
            .outp(out_6477)
        );        
        

        logic [WIDTH-1:0] out_6478;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6478 (
            .a(out_6476),
            .b(out_6477),
            .outp(out_6478)
        );        
        

        logic [WIDTH-1:0] out_6479;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6479 (
            .a(out_6470),
            .b(out_6478),
            .outp(out_6479)
        );        
        

        logic [WIDTH-1:0] out_6480;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.263484)
        ) inst_6480 (
            .outp(out_6480)
        );
        

        logic [WIDTH-1:0] out_6481;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6481 (
            .a(out_6480),
            .b(out_1826),
            .outp(out_6481)
        );        
        

        logic [WIDTH-1:0] out_6482;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6482 (
            .a(out_1823),
            .b(out_6481),
            .outp(out_6482)
        );        
        

        logic [WIDTH-1:0] out_6483;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.94178)
        ) inst_6483 (
            .outp(out_6483)
        );
        

        logic [WIDTH-1:0] out_6484;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6484 (
            .a(out_1831),
            .b(out_6483),
            .outp(out_6484)
        );        
        

        logic [WIDTH-1:0] out_6485;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6485 (
            .a(out_6482),
            .b(out_6484),
            .outp(out_6485)
        );        
        

        logic [WIDTH-1:0] out_6486;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.05264)
        ) inst_6486 (
            .outp(out_6486)
        );
        

        logic [WIDTH-1:0] out_6487;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6487 (
            .a(out_6486),
            .b(out_1834),
            .outp(out_6487)
        );        
        

        logic [WIDTH-1:0] out_6488;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6488 (
            .a(out_6485),
            .b(out_6487),
            .outp(out_6488)
        );        
        

        logic [WIDTH-1:0] out_6489;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6489 (
            .a(out_1834),
            .b(out_6486),
            .outp(out_6489)
        );        
        

        logic [WIDTH-1:0] out_6490;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6490 (
            .a(out_6483),
            .b(out_1831),
            .outp(out_6490)
        );        
        

        logic [WIDTH-1:0] out_6491;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6491 (
            .a(out_6489),
            .b(out_6490),
            .outp(out_6491)
        );        
        

        logic [WIDTH-1:0] out_6492;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6492 (
            .a(out_6481),
            .b(out_1823),
            .outp(out_6492)
        );        
        

        logic [WIDTH-1:0] out_6493;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6493 (
            .a(out_6491),
            .b(out_6492),
            .outp(out_6493)
        );        
        

        logic [WIDTH-1:0] out_6494;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6494 (
            .a(out_6488),
            .b(out_6493),
            .outp(out_6494)
        );        
        

        logic [WIDTH-1:0] out_6495;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6495 (
            .in(out_6494),
            .outp(out_6495)
        );
        

        logic [WIDTH-1:0] out_6496;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.075)
        ) inst_6496 (
            .outp(out_6496)
        );
        

        logic [WIDTH-1:0] out_6497;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6497 (
            .a(out_14),
            .b(out_6496),
            .outp(out_6497)
        );        
        

        logic [WIDTH-1:0] out_6498;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6498 (
            .in(out_6497),
            .outp(out_6498)
        );
        

        logic [WIDTH-1:0] out_6499;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.0255)
        ) inst_6499 (
            .outp(out_6499)
        );
        

        logic [WIDTH-1:0] out_6500;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6500 (
            .a(out_3),
            .b(out_6499),
            .outp(out_6500)
        );        
        

        logic [WIDTH-1:0] out_6501;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6501 (
            .in(out_6500),
            .outp(out_6501)
        );
        

        logic [WIDTH-1:0] out_6502;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6502 (
            .a(out_6498),
            .b(out_6501),
            .outp(out_6502)
        );        
        

        logic [WIDTH-1:0] out_6503;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6503 (
            .in(out_6502),
            .outp(out_6503)
        );
        

        logic [WIDTH-1:0] out_6504;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6504 (
            .a(out_9),
            .b(out_6503),
            .outp(out_6504)
        );        
        

        logic [WIDTH-1:0] out_6505;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6505 (
            .a(out_6495),
            .b(out_6504),
            .outp(out_6505)
        );        
        

        logic [WIDTH-1:0] out_6506;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6506 (
            .a(out_6503),
            .b(out_21),
            .outp(out_6506)
        );        
        

        logic [WIDTH-1:0] out_6507;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6507 (
            .a(out_6505),
            .b(out_6506),
            .outp(out_6507)
        );        
        

        logic [WIDTH-1:0] out_6508;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6508 (
            .a(out_6479),
            .b(out_6507),
            .outp(out_6508)
        );        
        

        logic [WIDTH-1:0] out_6509;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6509 (
            .a(out_14),
            .b(out_3253),
            .outp(out_6509)
        );        
        

        logic [WIDTH-1:0] out_6510;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6510 (
            .a(out_6462),
            .b(out_6509),
            .outp(out_6510)
        );        
        

        logic [WIDTH-1:0] out_6511;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.6255)
        ) inst_6511 (
            .outp(out_6511)
        );
        

        logic [WIDTH-1:0] out_6512;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6512 (
            .a(out_3),
            .b(out_6511),
            .outp(out_6512)
        );        
        

        logic [WIDTH-1:0] out_6513;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6513 (
            .a(out_6510),
            .b(out_6512),
            .outp(out_6513)
        );        
        

        logic [WIDTH-1:0] out_6514;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5255)
        ) inst_6514 (
            .outp(out_6514)
        );
        

        logic [WIDTH-1:0] out_6515;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6515 (
            .a(out_6514),
            .b(out_3),
            .outp(out_6515)
        );        
        

        logic [WIDTH-1:0] out_6516;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6516 (
            .a(out_6513),
            .b(out_6515),
            .outp(out_6516)
        );        
        

        logic [WIDTH-1:0] out_6517;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6517 (
            .a(out_6508),
            .b(out_6516),
            .outp(out_6517)
        );        
        

        logic [WIDTH-1:0] out_6518;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6518 (
            .a(out_14),
            .b(out_4157),
            .outp(out_6518)
        );        
        

        logic [WIDTH-1:0] out_6519;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6519 (
            .in(out_6518),
            .outp(out_6519)
        );
        

        logic [WIDTH-1:0] out_6520;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5755)
        ) inst_6520 (
            .outp(out_6520)
        );
        

        logic [WIDTH-1:0] out_6521;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6521 (
            .a(out_3),
            .b(out_6520),
            .outp(out_6521)
        );        
        

        logic [WIDTH-1:0] out_6522;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6522 (
            .in(out_6521),
            .outp(out_6522)
        );
        

        logic [WIDTH-1:0] out_6523;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6523 (
            .a(out_6519),
            .b(out_6522),
            .outp(out_6523)
        );        
        

        logic [WIDTH-1:0] out_6524;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6524 (
            .in(out_6523),
            .outp(out_6524)
        );
        

        logic [WIDTH-1:0] out_6525;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6525 (
            .a(out_6524),
            .b(out_460),
            .outp(out_6525)
        );        
        

        logic [WIDTH-1:0] out_6526;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6526 (
            .a(out_6517),
            .b(out_6525),
            .outp(out_6526)
        );        
        

        logic [WIDTH-1:0] out_6527;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6527 (
            .a(out_6215),
            .b(out_14),
            .outp(out_6527)
        );        
        

        logic [WIDTH-1:0] out_6528;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6528 (
            .a(out_6509),
            .b(out_6527),
            .outp(out_6528)
        );        
        

        logic [WIDTH-1:0] out_6529;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.4005)
        ) inst_6529 (
            .outp(out_6529)
        );
        

        logic [WIDTH-1:0] out_6530;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6530 (
            .a(out_3),
            .b(out_6529),
            .outp(out_6530)
        );        
        

        logic [WIDTH-1:0] out_6531;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6531 (
            .a(out_6528),
            .b(out_6530),
            .outp(out_6531)
        );        
        

        logic [WIDTH-1:0] out_6532;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.3005)
        ) inst_6532 (
            .outp(out_6532)
        );
        

        logic [WIDTH-1:0] out_6533;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6533 (
            .a(out_6532),
            .b(out_3),
            .outp(out_6533)
        );        
        

        logic [WIDTH-1:0] out_6534;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6534 (
            .a(out_6531),
            .b(out_6533),
            .outp(out_6534)
        );        
        

        logic [WIDTH-1:0] out_6535;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6535 (
            .a(out_6526),
            .b(out_6534),
            .outp(out_6535)
        );        
        

        logic [WIDTH-1:0] out_6536;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.1255)
        ) inst_6536 (
            .outp(out_6536)
        );
        

        logic [WIDTH-1:0] out_6537;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6537 (
            .a(out_3),
            .b(out_6536),
            .outp(out_6537)
        );        
        

        logic [WIDTH-1:0] out_6538;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6538 (
            .in(out_6537),
            .outp(out_6538)
        );
        

        logic [WIDTH-1:0] out_6539;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6539 (
            .a(out_6498),
            .b(out_6538),
            .outp(out_6539)
        );        
        

        logic [WIDTH-1:0] out_6540;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6540 (
            .in(out_6539),
            .outp(out_6540)
        );
        

        logic [WIDTH-1:0] out_6541;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6541 (
            .a(out_9),
            .b(out_6540),
            .outp(out_6541)
        );        
        

        logic [WIDTH-1:0] out_6542;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6542 (
            .a(out_6540),
            .b(out_21),
            .outp(out_6542)
        );        
        

        logic [WIDTH-1:0] out_6543;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6543 (
            .a(out_6541),
            .b(out_6542),
            .outp(out_6543)
        );        
        

        logic [WIDTH-1:0] out_6544;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6544 (
            .a(out_6535),
            .b(out_6543),
            .outp(out_6544)
        );        
        

        logic [WIDTH-1:0] out_6545;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.425)
        ) inst_6545 (
            .outp(out_6545)
        );
        

        logic [WIDTH-1:0] out_6546;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6546 (
            .a(out_6545),
            .b(out_14),
            .outp(out_6546)
        );        
        

        logic [WIDTH-1:0] out_6547;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6547 (
            .a(out_6530),
            .b(out_6546),
            .outp(out_6547)
        );        
        

        logic [WIDTH-1:0] out_6548;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.8505)
        ) inst_6548 (
            .outp(out_6548)
        );
        

        logic [WIDTH-1:0] out_6549;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6549 (
            .a(out_6548),
            .b(out_3),
            .outp(out_6549)
        );        
        

        logic [WIDTH-1:0] out_6550;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6550 (
            .a(out_6547),
            .b(out_6549),
            .outp(out_6550)
        );        
        

        logic [WIDTH-1:0] out_6551;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6551 (
            .in(out_6216),
            .outp(out_6551)
        );
        

        logic [WIDTH-1:0] out_6552;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6552 (
            .a(out_6538),
            .b(out_6551),
            .outp(out_6552)
        );        
        

        logic [WIDTH-1:0] out_6553;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6553 (
            .in(out_6552),
            .outp(out_6553)
        );
        

        logic [WIDTH-1:0] out_6554;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6554 (
            .a(out_9),
            .b(out_6553),
            .outp(out_6554)
        );        
        

        logic [WIDTH-1:0] out_6555;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6555 (
            .a(out_6550),
            .b(out_6554),
            .outp(out_6555)
        );        
        

        logic [WIDTH-1:0] out_6556;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6556 (
            .a(out_6553),
            .b(out_21),
            .outp(out_6556)
        );        
        

        logic [WIDTH-1:0] out_6557;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6557 (
            .a(out_6555),
            .b(out_6556),
            .outp(out_6557)
        );        
        

        logic [WIDTH-1:0] out_6558;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6558 (
            .a(out_6557),
            .b(out_6216),
            .outp(out_6558)
        );        
        

        logic [WIDTH-1:0] out_6559;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6559 (
            .a(out_6544),
            .b(out_6558),
            .outp(out_6559)
        );        
        

        logic [WIDTH-1:0] out_6560;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.242)
        ) inst_6560 (
            .outp(out_6560)
        );
        

        logic [WIDTH-1:0] out_6561;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6561 (
            .a(out_6560),
            .b(out_3),
            .outp(out_6561)
        );        
        

        logic [WIDTH-1:0] out_6562;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.742)
        ) inst_6562 (
            .outp(out_6562)
        );
        

        logic [WIDTH-1:0] out_6563;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6563 (
            .a(out_6562),
            .b(out_3),
            .outp(out_6563)
        );        
        

        logic [WIDTH-1:0] out_6564;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6564 (
            .in(out_6563),
            .outp(out_6564)
        );
        

        logic [WIDTH-1:0] out_6565;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6565 (
            .a(out_6561),
            .b(out_6564),
            .outp(out_6565)
        );        
        

        logic [WIDTH-1:0] out_6566;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6566 (
            .a(out_6565),
            .b(out_6343),
            .outp(out_6566)
        );        
        

        logic [WIDTH-1:0] out_6567;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6567 (
            .a(out_6566),
            .b(out_6345),
            .outp(out_6567)
        );        
        

        logic [WIDTH-1:0] out_6568;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.517)
        ) inst_6568 (
            .outp(out_6568)
        );
        

        logic [WIDTH-1:0] out_6569;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6569 (
            .a(out_6568),
            .b(out_3),
            .outp(out_6569)
        );        
        

        logic [WIDTH-1:0] out_6570;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6570 (
            .in(out_6569),
            .outp(out_6570)
        );
        

        logic [WIDTH-1:0] out_6571;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6571 (
            .a(out_6570),
            .b(out_6061),
            .outp(out_6571)
        );        
        

        logic [WIDTH-1:0] out_6572;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6572 (
            .in(out_6571),
            .outp(out_6572)
        );
        

        logic [WIDTH-1:0] out_6573;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6573 (
            .a(out_6572),
            .b(out_21),
            .outp(out_6573)
        );        
        

        logic [WIDTH-1:0] out_6574;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.8578)
        ) inst_6574 (
            .outp(out_6574)
        );
        

        logic [WIDTH-1:0] out_6575;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6575 (
            .a(out_6574),
            .b(out_556),
            .outp(out_6575)
        );        
        

        logic [WIDTH-1:0] out_6576;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6576 (
            .a(out_6575),
            .b(out_559),
            .outp(out_6576)
        );        
        

        logic [WIDTH-1:0] out_6577;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.1972)
        ) inst_6577 (
            .outp(out_6577)
        );
        

        logic [WIDTH-1:0] out_6578;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6578 (
            .a(out_6577),
            .b(out_2653),
            .outp(out_6578)
        );        
        

        logic [WIDTH-1:0] out_6579;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6579 (
            .a(out_6576),
            .b(out_6578),
            .outp(out_6579)
        );        
        

        logic [WIDTH-1:0] out_6580;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6580 (
            .a(out_6579),
            .b(out_6360),
            .outp(out_6580)
        );        
        

        logic [WIDTH-1:0] out_6581;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6581 (
            .a(out_2653),
            .b(out_6577),
            .outp(out_6581)
        );        
        

        logic [WIDTH-1:0] out_6582;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6582 (
            .a(out_559),
            .b(out_6575),
            .outp(out_6582)
        );        
        

        logic [WIDTH-1:0] out_6583;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6583 (
            .a(out_6581),
            .b(out_6582),
            .outp(out_6583)
        );        
        

        logic [WIDTH-1:0] out_6584;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6584 (
            .a(out_6583),
            .b(out_6365),
            .outp(out_6584)
        );        
        

        logic [WIDTH-1:0] out_6585;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6585 (
            .a(out_6580),
            .b(out_6584),
            .outp(out_6585)
        );        
        

        logic [WIDTH-1:0] out_6586;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6586 (
            .in(out_6585),
            .outp(out_6586)
        );
        

        logic [WIDTH-1:0] out_6587;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6587 (
            .a(out_6573),
            .b(out_6586),
            .outp(out_6587)
        );        
        

        logic [WIDTH-1:0] out_6588;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6588 (
            .a(out_9),
            .b(out_6572),
            .outp(out_6588)
        );        
        

        logic [WIDTH-1:0] out_6589;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6589 (
            .a(out_6587),
            .b(out_6588),
            .outp(out_6589)
        );        
        

        logic [WIDTH-1:0] out_6590;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6590 (
            .a(out_6567),
            .b(out_6589),
            .outp(out_6590)
        );        
        

        logic [WIDTH-1:0] out_6591;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6591 (
            .a(out_6573),
            .b(out_6590),
            .outp(out_6591)
        );        
        

        logic [WIDTH-1:0] out_6592;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6592 (
            .a(out_6559),
            .b(out_6591),
            .outp(out_6592)
        );        
        

        logic [WIDTH-1:0] out_6593;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.15)
        ) inst_6593 (
            .outp(out_6593)
        );
        

        logic [WIDTH-1:0] out_6594;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6594 (
            .a(out_6593),
            .b(out_3),
            .outp(out_6594)
        );        
        

        logic [WIDTH-1:0] out_6595;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6595 (
            .a(out_6073),
            .b(out_3),
            .outp(out_6595)
        );        
        

        logic [WIDTH-1:0] out_6596;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6596 (
            .in(out_6595),
            .outp(out_6596)
        );
        

        logic [WIDTH-1:0] out_6597;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6597 (
            .a(out_6594),
            .b(out_6596),
            .outp(out_6597)
        );        
        

        logic [WIDTH-1:0] out_6598;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6598 (
            .a(out_6597),
            .b(out_6088),
            .outp(out_6598)
        );        
        

        logic [WIDTH-1:0] out_6599;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6599 (
            .a(out_6598),
            .b(out_6074),
            .outp(out_6599)
        );        
        

        logic [WIDTH-1:0] out_6600;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6600 (
            .a(out_6592),
            .b(out_6599),
            .outp(out_6600)
        );        
        

        logic [WIDTH-1:0] out_6601;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.95)
        ) inst_6601 (
            .outp(out_6601)
        );
        

        logic [WIDTH-1:0] out_6602;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6602 (
            .a(out_6601),
            .b(out_194),
            .outp(out_6602)
        );        
        

        logic [WIDTH-1:0] out_6603;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.5)
        ) inst_6603 (
            .outp(out_6603)
        );
        

        logic [WIDTH-1:0] out_6604;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6604 (
            .a(out_6603),
            .b(out_194),
            .outp(out_6604)
        );        
        

        logic [WIDTH-1:0] out_6605;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6605 (
            .in(out_6604),
            .outp(out_6605)
        );
        

        logic [WIDTH-1:0] out_6606;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6606 (
            .a(out_6602),
            .b(out_6605),
            .outp(out_6606)
        );        
        

        logic [WIDTH-1:0] out_6607;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.6875)
        ) inst_6607 (
            .outp(out_6607)
        );
        

        logic [WIDTH-1:0] out_6608;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6608 (
            .a(out_6607),
            .b(out_204),
            .outp(out_6608)
        );        
        

        logic [WIDTH-1:0] out_6609;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6609 (
            .in(out_6608),
            .outp(out_6609)
        );
        

        logic [WIDTH-1:0] out_6610;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6610 (
            .a(out_6391),
            .b(out_6609),
            .outp(out_6610)
        );        
        

        logic [WIDTH-1:0] out_6611;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6611 (
            .in(out_6610),
            .outp(out_6611)
        );
        

        logic [WIDTH-1:0] out_6612;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6612 (
            .a(out_200),
            .b(out_6611),
            .outp(out_6612)
        );        
        

        logic [WIDTH-1:0] out_6613;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6613 (
            .a(out_6606),
            .b(out_6612),
            .outp(out_6613)
        );        
        

        logic [WIDTH-1:0] out_6614;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6614 (
            .in(out_6602),
            .outp(out_6614)
        );
        

        logic [WIDTH-1:0] out_6615;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6615 (
            .a(out_6391),
            .b(out_6614),
            .outp(out_6615)
        );        
        

        logic [WIDTH-1:0] out_6616;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6616 (
            .in(out_6615),
            .outp(out_6616)
        );
        

        logic [WIDTH-1:0] out_6617;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6617 (
            .a(out_6616),
            .b(out_214),
            .outp(out_6617)
        );        
        

        logic [WIDTH-1:0] out_6618;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6618 (
            .a(out_6613),
            .b(out_6617),
            .outp(out_6618)
        );        
        

        logic [WIDTH-1:0] out_6619;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6619 (
            .a(out_6618),
            .b(out_6088),
            .outp(out_6619)
        );        
        

        logic [WIDTH-1:0] out_6620;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6620 (
            .a(out_6619),
            .b(out_6074),
            .outp(out_6620)
        );        
        

        logic [WIDTH-1:0] out_6621;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6621 (
            .a(out_6600),
            .b(out_6620),
            .outp(out_6621)
        );        
        

        logic [WIDTH-1:0] out_6622;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.35)
        ) inst_6622 (
            .outp(out_6622)
        );
        

        logic [WIDTH-1:0] out_6623;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6623 (
            .a(out_6622),
            .b(out_3),
            .outp(out_6623)
        );        
        

        logic [WIDTH-1:0] out_6624;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.85)
        ) inst_6624 (
            .outp(out_6624)
        );
        

        logic [WIDTH-1:0] out_6625;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6625 (
            .a(out_6624),
            .b(out_3),
            .outp(out_6625)
        );        
        

        logic [WIDTH-1:0] out_6626;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6626 (
            .in(out_6625),
            .outp(out_6626)
        );
        

        logic [WIDTH-1:0] out_6627;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6627 (
            .a(out_6623),
            .b(out_6626),
            .outp(out_6627)
        );        
        

        logic [WIDTH-1:0] out_6628;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6628 (
            .a(out_6627),
            .b(out_6343),
            .outp(out_6628)
        );        
        

        logic [WIDTH-1:0] out_6629;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6629 (
            .a(out_6628),
            .b(out_6345),
            .outp(out_6629)
        );        
        

        logic [WIDTH-1:0] out_6630;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.625)
        ) inst_6630 (
            .outp(out_6630)
        );
        

        logic [WIDTH-1:0] out_6631;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6631 (
            .a(out_6630),
            .b(out_3),
            .outp(out_6631)
        );        
        

        logic [WIDTH-1:0] out_6632;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6632 (
            .in(out_6631),
            .outp(out_6632)
        );
        

        logic [WIDTH-1:0] out_6633;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6633 (
            .a(out_6632),
            .b(out_6061),
            .outp(out_6633)
        );        
        

        logic [WIDTH-1:0] out_6634;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6634 (
            .in(out_6633),
            .outp(out_6634)
        );
        

        logic [WIDTH-1:0] out_6635;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6635 (
            .a(out_6634),
            .b(out_21),
            .outp(out_6635)
        );        
        

        logic [WIDTH-1:0] out_6636;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.1625)
        ) inst_6636 (
            .outp(out_6636)
        );
        

        logic [WIDTH-1:0] out_6637;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6637 (
            .a(out_6636),
            .b(out_556),
            .outp(out_6637)
        );        
        

        logic [WIDTH-1:0] out_6638;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6638 (
            .a(out_6637),
            .b(out_559),
            .outp(out_6638)
        );        
        

        logic [WIDTH-1:0] out_6639;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.8925)
        ) inst_6639 (
            .outp(out_6639)
        );
        

        logic [WIDTH-1:0] out_6640;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6640 (
            .a(out_6639),
            .b(out_2653),
            .outp(out_6640)
        );        
        

        logic [WIDTH-1:0] out_6641;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6641 (
            .a(out_6638),
            .b(out_6640),
            .outp(out_6641)
        );        
        

        logic [WIDTH-1:0] out_6642;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6642 (
            .a(out_6641),
            .b(out_6360),
            .outp(out_6642)
        );        
        

        logic [WIDTH-1:0] out_6643;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6643 (
            .a(out_2653),
            .b(out_6639),
            .outp(out_6643)
        );        
        

        logic [WIDTH-1:0] out_6644;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6644 (
            .a(out_559),
            .b(out_6637),
            .outp(out_6644)
        );        
        

        logic [WIDTH-1:0] out_6645;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6645 (
            .a(out_6643),
            .b(out_6644),
            .outp(out_6645)
        );        
        

        logic [WIDTH-1:0] out_6646;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6646 (
            .a(out_6645),
            .b(out_6365),
            .outp(out_6646)
        );        
        

        logic [WIDTH-1:0] out_6647;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6647 (
            .a(out_6642),
            .b(out_6646),
            .outp(out_6647)
        );        
        

        logic [WIDTH-1:0] out_6648;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6648 (
            .in(out_6647),
            .outp(out_6648)
        );
        

        logic [WIDTH-1:0] out_6649;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6649 (
            .a(out_6635),
            .b(out_6648),
            .outp(out_6649)
        );        
        

        logic [WIDTH-1:0] out_6650;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6650 (
            .a(out_9),
            .b(out_6634),
            .outp(out_6650)
        );        
        

        logic [WIDTH-1:0] out_6651;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6651 (
            .a(out_6649),
            .b(out_6650),
            .outp(out_6651)
        );        
        

        logic [WIDTH-1:0] out_6652;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6652 (
            .a(out_6629),
            .b(out_6651),
            .outp(out_6652)
        );        
        

        logic [WIDTH-1:0] out_6653;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6653 (
            .a(out_6635),
            .b(out_6652),
            .outp(out_6653)
        );        
        

        logic [WIDTH-1:0] out_6654;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6654 (
            .a(out_6621),
            .b(out_6653),
            .outp(out_6654)
        );        
        

        logic [WIDTH-1:0] out_6655;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.05)
        ) inst_6655 (
            .outp(out_6655)
        );
        

        logic [WIDTH-1:0] out_6656;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6656 (
            .a(out_6655),
            .b(out_3),
            .outp(out_6656)
        );        
        

        logic [WIDTH-1:0] out_6657;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.15)
        ) inst_6657 (
            .outp(out_6657)
        );
        

        logic [WIDTH-1:0] out_6658;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6658 (
            .a(out_6657),
            .b(out_3),
            .outp(out_6658)
        );        
        

        logic [WIDTH-1:0] out_6659;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6659 (
            .in(out_6658),
            .outp(out_6659)
        );
        

        logic [WIDTH-1:0] out_6660;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6660 (
            .a(out_6656),
            .b(out_6659),
            .outp(out_6660)
        );        
        

        logic [WIDTH-1:0] out_6661;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6661 (
            .a(out_6660),
            .b(out_6088),
            .outp(out_6661)
        );        
        

        logic [WIDTH-1:0] out_6662;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6662 (
            .a(out_6661),
            .b(out_6060),
            .outp(out_6662)
        );        
        

        logic [WIDTH-1:0] out_6663;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6663 (
            .a(out_6654),
            .b(out_6662),
            .outp(out_6663)
        );        
        

        logic [WIDTH-1:0] out_6664;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6664 (
            .a(out_4158),
            .b(out_4162),
            .outp(out_6664)
        );        
        

        logic [WIDTH-1:0] out_6665;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6665 (
            .a(out_6664),
            .b(out_6216),
            .outp(out_6665)
        );        
        

        logic [WIDTH-1:0] out_6666;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6666 (
            .a(out_6665),
            .b(out_6088),
            .outp(out_6666)
        );        
        

        logic [WIDTH-1:0] out_6667;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6667 (
            .a(out_6663),
            .b(out_6666),
            .outp(out_6667)
        );        
        

        logic [WIDTH-1:0] out_6668;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6668 (
            .a(out_4162),
            .b(out_6656),
            .outp(out_6668)
        );        
        

        logic [WIDTH-1:0] out_6669;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6669 (
            .a(out_1851),
            .b(out_6061),
            .outp(out_6669)
        );        
        

        logic [WIDTH-1:0] out_6670;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6670 (
            .in(out_6669),
            .outp(out_6670)
        );
        

        logic [WIDTH-1:0] out_6671;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6671 (
            .a(out_9),
            .b(out_6670),
            .outp(out_6671)
        );        
        

        logic [WIDTH-1:0] out_6672;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6672 (
            .a(out_6668),
            .b(out_6671),
            .outp(out_6672)
        );        
        

        logic [WIDTH-1:0] out_6673;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6673 (
            .a(out_6670),
            .b(out_21),
            .outp(out_6673)
        );        
        

        logic [WIDTH-1:0] out_6674;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6674 (
            .a(out_6672),
            .b(out_6673),
            .outp(out_6674)
        );        
        

        logic [WIDTH-1:0] out_6675;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6675 (
            .a(out_6674),
            .b(out_6422),
            .outp(out_6675)
        );        
        

        logic [WIDTH-1:0] out_6676;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6676 (
            .a(out_6675),
            .b(out_6074),
            .outp(out_6676)
        );        
        

        logic [WIDTH-1:0] out_6677;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6677 (
            .a(out_6667),
            .b(out_6676),
            .outp(out_6677)
        );        
        

        logic [WIDTH-1:0] out_6678;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.7)
        ) inst_6678 (
            .outp(out_6678)
        );
        

        logic [WIDTH-1:0] out_6679;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6679 (
            .a(out_6678),
            .b(out_14),
            .outp(out_6679)
        );        
        

        logic [WIDTH-1:0] out_6680;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6680 (
            .a(out_6477),
            .b(out_6679),
            .outp(out_6680)
        );        
        

        logic [WIDTH-1:0] out_6681;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6681 (
            .a(out_6680),
            .b(out_6465),
            .outp(out_6681)
        );        
        

        logic [WIDTH-1:0] out_6682;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6682 (
            .a(out_6681),
            .b(out_6468),
            .outp(out_6682)
        );        
        

        logic [WIDTH-1:0] out_6683;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6683 (
            .a(out_6677),
            .b(out_6682),
            .outp(out_6683)
        );        
        

        logic [WIDTH-1:0] out_6684;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.9705)
        ) inst_6684 (
            .outp(out_6684)
        );
        

        logic [WIDTH-1:0] out_6685;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6685 (
            .a(out_3),
            .b(out_6684),
            .outp(out_6685)
        );        
        

        logic [WIDTH-1:0] out_6686;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6686 (
            .a(out_6528),
            .b(out_6685),
            .outp(out_6686)
        );        
        

        logic [WIDTH-1:0] out_6687;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.8705)
        ) inst_6687 (
            .outp(out_6687)
        );
        

        logic [WIDTH-1:0] out_6688;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6688 (
            .a(out_6687),
            .b(out_3),
            .outp(out_6688)
        );        
        

        logic [WIDTH-1:0] out_6689;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6689 (
            .a(out_6686),
            .b(out_6688),
            .outp(out_6689)
        );        
        

        logic [WIDTH-1:0] out_6690;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6690 (
            .a(out_6683),
            .b(out_6689),
            .outp(out_6690)
        );        
        

        logic [WIDTH-1:0] out_6691;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.695499)
        ) inst_6691 (
            .outp(out_6691)
        );
        

        logic [WIDTH-1:0] out_6692;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6692 (
            .a(out_3),
            .b(out_6691),
            .outp(out_6692)
        );        
        

        logic [WIDTH-1:0] out_6693;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6693 (
            .in(out_6692),
            .outp(out_6693)
        );
        

        logic [WIDTH-1:0] out_6694;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6694 (
            .a(out_6498),
            .b(out_6693),
            .outp(out_6694)
        );        
        

        logic [WIDTH-1:0] out_6695;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6695 (
            .in(out_6694),
            .outp(out_6695)
        );
        

        logic [WIDTH-1:0] out_6696;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6696 (
            .a(out_9),
            .b(out_6695),
            .outp(out_6696)
        );        
        

        logic [WIDTH-1:0] out_6697;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6697 (
            .a(out_6695),
            .b(out_21),
            .outp(out_6697)
        );        
        

        logic [WIDTH-1:0] out_6698;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6698 (
            .a(out_6696),
            .b(out_6697),
            .outp(out_6698)
        );        
        

        logic [WIDTH-1:0] out_6699;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6699 (
            .a(out_6690),
            .b(out_6698),
            .outp(out_6699)
        );        
        

        logic [WIDTH-1:0] out_6700;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6700 (
            .a(out_6546),
            .b(out_6685),
            .outp(out_6700)
        );        
        

        logic [WIDTH-1:0] out_6701;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.4205)
        ) inst_6701 (
            .outp(out_6701)
        );
        

        logic [WIDTH-1:0] out_6702;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6702 (
            .a(out_6701),
            .b(out_3),
            .outp(out_6702)
        );        
        

        logic [WIDTH-1:0] out_6703;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6703 (
            .a(out_6700),
            .b(out_6702),
            .outp(out_6703)
        );        
        

        logic [WIDTH-1:0] out_6704;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6704 (
            .a(out_6551),
            .b(out_6693),
            .outp(out_6704)
        );        
        

        logic [WIDTH-1:0] out_6705;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6705 (
            .in(out_6704),
            .outp(out_6705)
        );
        

        logic [WIDTH-1:0] out_6706;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6706 (
            .a(out_9),
            .b(out_6705),
            .outp(out_6706)
        );        
        

        logic [WIDTH-1:0] out_6707;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6707 (
            .a(out_6703),
            .b(out_6706),
            .outp(out_6707)
        );        
        

        logic [WIDTH-1:0] out_6708;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6708 (
            .a(out_6705),
            .b(out_21),
            .outp(out_6708)
        );        
        

        logic [WIDTH-1:0] out_6709;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6709 (
            .a(out_6707),
            .b(out_6708),
            .outp(out_6709)
        );        
        

        logic [WIDTH-1:0] out_6710;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6710 (
            .a(out_6709),
            .b(out_6216),
            .outp(out_6710)
        );        
        

        logic [WIDTH-1:0] out_6711;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6711 (
            .a(out_6699),
            .b(out_6710),
            .outp(out_6711)
        );        
        

        logic [WIDTH-1:0] out_6712;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.320499)
        ) inst_6712 (
            .outp(out_6712)
        );
        

        logic [WIDTH-1:0] out_6713;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6713 (
            .a(out_3),
            .b(out_6712),
            .outp(out_6713)
        );        
        

        logic [WIDTH-1:0] out_6714;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6714 (
            .a(out_6510),
            .b(out_6713),
            .outp(out_6714)
        );        
        

        logic [WIDTH-1:0] out_6715;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.220499)
        ) inst_6715 (
            .outp(out_6715)
        );
        

        logic [WIDTH-1:0] out_6716;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6716 (
            .a(out_6715),
            .b(out_3),
            .outp(out_6716)
        );        
        

        logic [WIDTH-1:0] out_6717;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6717 (
            .a(out_6714),
            .b(out_6716),
            .outp(out_6717)
        );        
        

        logic [WIDTH-1:0] out_6718;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6718 (
            .a(out_6711),
            .b(out_6717),
            .outp(out_6718)
        );        
        

        logic [WIDTH-1:0] out_6719;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.129501)
        ) inst_6719 (
            .outp(out_6719)
        );
        

        logic [WIDTH-1:0] out_6720;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6720 (
            .a(out_6719),
            .b(out_3),
            .outp(out_6720)
        );        
        

        logic [WIDTH-1:0] out_6721;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6721 (
            .a(out_6509),
            .b(out_6720),
            .outp(out_6721)
        );        
        

        logic [WIDTH-1:0] out_6722;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.229501)
        ) inst_6722 (
            .outp(out_6722)
        );
        

        logic [WIDTH-1:0] out_6723;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6723 (
            .a(out_6722),
            .b(out_3),
            .outp(out_6723)
        );        
        

        logic [WIDTH-1:0] out_6724;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6724 (
            .in(out_6723),
            .outp(out_6724)
        );
        

        logic [WIDTH-1:0] out_6725;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6725 (
            .a(out_6721),
            .b(out_6724),
            .outp(out_6725)
        );        
        

        logic [WIDTH-1:0] out_6726;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6726 (
            .a(out_6496),
            .b(out_14),
            .outp(out_6726)
        );        
        

        logic [WIDTH-1:0] out_6727;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6727 (
            .a(out_6725),
            .b(out_6726),
            .outp(out_6727)
        );        
        

        logic [WIDTH-1:0] out_6728;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6728 (
            .a(out_6718),
            .b(out_6727),
            .outp(out_6728)
        );        
        

        logic [WIDTH-1:0] out_6729;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6729 (
            .a(out_6462),
            .b(out_6497),
            .outp(out_6729)
        );        
        

        logic [WIDTH-1:0] out_6730;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6730 (
            .a(out_6729),
            .b(out_6713),
            .outp(out_6730)
        );        
        

        logic [WIDTH-1:0] out_6731;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6731 (
            .a(out_6730),
            .b(out_6724),
            .outp(out_6731)
        );        
        

        logic [WIDTH-1:0] out_6732;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.0454988)
        ) inst_6732 (
            .outp(out_6732)
        );
        

        logic [WIDTH-1:0] out_6733;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6733 (
            .a(out_3),
            .b(out_6732),
            .outp(out_6733)
        );        
        

        logic [WIDTH-1:0] out_6734;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6734 (
            .in(out_6733),
            .outp(out_6734)
        );
        

        logic [WIDTH-1:0] out_6735;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6735 (
            .a(out_6498),
            .b(out_6734),
            .outp(out_6735)
        );        
        

        logic [WIDTH-1:0] out_6736;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6736 (
            .in(out_6735),
            .outp(out_6736)
        );
        

        logic [WIDTH-1:0] out_6737;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6737 (
            .a(out_9),
            .b(out_6736),
            .outp(out_6737)
        );        
        

        logic [WIDTH-1:0] out_6738;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6738 (
            .a(out_6731),
            .b(out_6737),
            .outp(out_6738)
        );        
        

        logic [WIDTH-1:0] out_6739;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6739 (
            .a(out_6736),
            .b(out_21),
            .outp(out_6739)
        );        
        

        logic [WIDTH-1:0] out_6740;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6740 (
            .a(out_6738),
            .b(out_6739),
            .outp(out_6740)
        );        
        

        logic [WIDTH-1:0] out_6741;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6741 (
            .a(out_6728),
            .b(out_6740),
            .outp(out_6741)
        );        
        

        logic [WIDTH-1:0] out_6742;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.604501)
        ) inst_6742 (
            .outp(out_6742)
        );
        

        logic [WIDTH-1:0] out_6743;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6743 (
            .a(out_6742),
            .b(out_3),
            .outp(out_6743)
        );        
        

        logic [WIDTH-1:0] out_6744;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6744 (
            .in(out_6743),
            .outp(out_6744)
        );
        

        logic [WIDTH-1:0] out_6745;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6745 (
            .a(out_6498),
            .b(out_6744),
            .outp(out_6745)
        );        
        

        logic [WIDTH-1:0] out_6746;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6746 (
            .in(out_6745),
            .outp(out_6746)
        );
        

        logic [WIDTH-1:0] out_6747;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6747 (
            .a(out_9),
            .b(out_6746),
            .outp(out_6747)
        );        
        

        logic [WIDTH-1:0] out_6748;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6748 (
            .a(out_6746),
            .b(out_21),
            .outp(out_6748)
        );        
        

        logic [WIDTH-1:0] out_6749;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6749 (
            .a(out_6747),
            .b(out_6748),
            .outp(out_6749)
        );        
        

        logic [WIDTH-1:0] out_6750;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6750 (
            .a(out_6741),
            .b(out_6749),
            .outp(out_6750)
        );        
        

        logic [WIDTH-1:0] out_6751;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.2375)
        ) inst_6751 (
            .outp(out_6751)
        );
        

        logic [WIDTH-1:0] out_6752;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6752 (
            .a(out_6751),
            .b(out_3),
            .outp(out_6752)
        );        
        

        logic [WIDTH-1:0] out_6753;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6753 (
            .a(out_6510),
            .b(out_6752),
            .outp(out_6753)
        );        
        

        logic [WIDTH-1:0] out_6754;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.3375)
        ) inst_6754 (
            .outp(out_6754)
        );
        

        logic [WIDTH-1:0] out_6755;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6755 (
            .a(out_6754),
            .b(out_3),
            .outp(out_6755)
        );        
        

        logic [WIDTH-1:0] out_6756;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6756 (
            .in(out_6755),
            .outp(out_6756)
        );
        

        logic [WIDTH-1:0] out_6757;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6757 (
            .a(out_6753),
            .b(out_6756),
            .outp(out_6757)
        );        
        

        logic [WIDTH-1:0] out_6758;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6758 (
            .a(out_6750),
            .b(out_6757),
            .outp(out_6758)
        );        
        

        logic [WIDTH-1:0] out_6759;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.36071)
        ) inst_6759 (
            .outp(out_6759)
        );
        

        logic [WIDTH-1:0] out_6760;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6760 (
            .a(out_6759),
            .b(out_194),
            .outp(out_6760)
        );        
        

        logic [WIDTH-1:0] out_6761;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6761 (
            .a(out_6510),
            .b(out_6760),
            .outp(out_6761)
        );        
        

        logic [WIDTH-1:0] out_6762;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.91072)
        ) inst_6762 (
            .outp(out_6762)
        );
        

        logic [WIDTH-1:0] out_6763;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6763 (
            .a(out_6762),
            .b(out_194),
            .outp(out_6763)
        );        
        

        logic [WIDTH-1:0] out_6764;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6764 (
            .in(out_6763),
            .outp(out_6764)
        );
        

        logic [WIDTH-1:0] out_6765;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6765 (
            .a(out_6761),
            .b(out_6764),
            .outp(out_6765)
        );        
        

        logic [WIDTH-1:0] out_6766;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6766 (
            .a(out_14),
            .b(out_6461),
            .outp(out_6766)
        );        
        

        logic [WIDTH-1:0] out_6767;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6767 (
            .in(out_6766),
            .outp(out_6767)
        );
        

        logic [WIDTH-1:0] out_6768;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.70089)
        ) inst_6768 (
            .outp(out_6768)
        );
        

        logic [WIDTH-1:0] out_6769;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6769 (
            .a(out_6768),
            .b(out_204),
            .outp(out_6769)
        );        
        

        logic [WIDTH-1:0] out_6770;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6770 (
            .in(out_6769),
            .outp(out_6770)
        );
        

        logic [WIDTH-1:0] out_6771;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6771 (
            .a(out_6767),
            .b(out_6770),
            .outp(out_6771)
        );        
        

        logic [WIDTH-1:0] out_6772;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6772 (
            .in(out_6771),
            .outp(out_6772)
        );
        

        logic [WIDTH-1:0] out_6773;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6773 (
            .a(out_200),
            .b(out_6772),
            .outp(out_6773)
        );        
        

        logic [WIDTH-1:0] out_6774;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6774 (
            .a(out_6765),
            .b(out_6773),
            .outp(out_6774)
        );        
        

        logic [WIDTH-1:0] out_6775;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6775 (
            .in(out_6760),
            .outp(out_6775)
        );
        

        logic [WIDTH-1:0] out_6776;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6776 (
            .a(out_6767),
            .b(out_6775),
            .outp(out_6776)
        );        
        

        logic [WIDTH-1:0] out_6777;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6777 (
            .in(out_6776),
            .outp(out_6777)
        );
        

        logic [WIDTH-1:0] out_6778;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6778 (
            .a(out_6777),
            .b(out_214),
            .outp(out_6778)
        );        
        

        logic [WIDTH-1:0] out_6779;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6779 (
            .a(out_6774),
            .b(out_6778),
            .outp(out_6779)
        );        
        

        logic [WIDTH-1:0] out_6780;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6780 (
            .a(out_6758),
            .b(out_6779),
            .outp(out_6780)
        );        
        

        logic [WIDTH-1:0] out_6781;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6781 (
            .a(out_14),
            .b(out_6657),
            .outp(out_6781)
        );        
        

        logic [WIDTH-1:0] out_6782;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6782 (
            .a(out_6462),
            .b(out_6781),
            .outp(out_6782)
        );        
        

        logic [WIDTH-1:0] out_6783;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.7305)
        ) inst_6783 (
            .outp(out_6783)
        );
        

        logic [WIDTH-1:0] out_6784;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6784 (
            .a(out_3),
            .b(out_6783),
            .outp(out_6784)
        );        
        

        logic [WIDTH-1:0] out_6785;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6785 (
            .a(out_6782),
            .b(out_6784),
            .outp(out_6785)
        );        
        

        logic [WIDTH-1:0] out_6786;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6305)
        ) inst_6786 (
            .outp(out_6786)
        );
        

        logic [WIDTH-1:0] out_6787;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6787 (
            .a(out_6786),
            .b(out_3),
            .outp(out_6787)
        );        
        

        logic [WIDTH-1:0] out_6788;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6788 (
            .a(out_6785),
            .b(out_6787),
            .outp(out_6788)
        );        
        

        logic [WIDTH-1:0] out_6789;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6789 (
            .a(out_6780),
            .b(out_6788),
            .outp(out_6789)
        );        
        

        logic [WIDTH-1:0] out_6790;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.71336)
        ) inst_6790 (
            .outp(out_6790)
        );
        

        logic [WIDTH-1:0] out_6791;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6791 (
            .a(out_6790),
            .b(out_1495),
            .outp(out_6791)
        );        
        

        logic [WIDTH-1:0] out_6792;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6792 (
            .a(out_3),
            .b(out_6791),
            .outp(out_6792)
        );        
        

        logic [WIDTH-1:0] out_6793;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6793 (
            .in(out_6792),
            .outp(out_6793)
        );
        

        logic [WIDTH-1:0] out_6794;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6794 (
            .a(out_6498),
            .b(out_6793),
            .outp(out_6794)
        );        
        

        logic [WIDTH-1:0] out_6795;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6795 (
            .in(out_6794),
            .outp(out_6795)
        );
        

        logic [WIDTH-1:0] out_6796;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6796 (
            .a(out_9),
            .b(out_6795),
            .outp(out_6796)
        );        
        

        logic [WIDTH-1:0] out_6797;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6797 (
            .a(out_6795),
            .b(out_21),
            .outp(out_6797)
        );        
        

        logic [WIDTH-1:0] out_6798;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6798 (
            .a(out_6796),
            .b(out_6797),
            .outp(out_6798)
        );        
        

        logic [WIDTH-1:0] out_6799;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6799 (
            .a(out_6789),
            .b(out_6798),
            .outp(out_6799)
        );        
        

        logic [WIDTH-1:0] out_6800;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.0705)
        ) inst_6800 (
            .outp(out_6800)
        );
        

        logic [WIDTH-1:0] out_6801;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6801 (
            .a(out_3),
            .b(out_6800),
            .outp(out_6801)
        );        
        

        logic [WIDTH-1:0] out_6802;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6802 (
            .a(out_6782),
            .b(out_6801),
            .outp(out_6802)
        );        
        

        logic [WIDTH-1:0] out_6803;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6803 (
            .a(out_3565),
            .b(out_3),
            .outp(out_6803)
        );        
        

        logic [WIDTH-1:0] out_6804;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6804 (
            .a(out_6802),
            .b(out_6803),
            .outp(out_6804)
        );        
        

        logic [WIDTH-1:0] out_6805;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6805 (
            .a(out_6799),
            .b(out_6804),
            .outp(out_6805)
        );        
        

        logic [WIDTH-1:0] out_6806;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8205)
        ) inst_6806 (
            .outp(out_6806)
        );
        

        logic [WIDTH-1:0] out_6807;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6807 (
            .a(out_3),
            .b(out_6806),
            .outp(out_6807)
        );        
        

        logic [WIDTH-1:0] out_6808;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6808 (
            .a(out_6782),
            .b(out_6807),
            .outp(out_6808)
        );        
        

        logic [WIDTH-1:0] out_6809;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.7205)
        ) inst_6809 (
            .outp(out_6809)
        );
        

        logic [WIDTH-1:0] out_6810;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6810 (
            .a(out_6809),
            .b(out_3),
            .outp(out_6810)
        );        
        

        logic [WIDTH-1:0] out_6811;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6811 (
            .a(out_6808),
            .b(out_6810),
            .outp(out_6811)
        );        
        

        logic [WIDTH-1:0] out_6812;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6812 (
            .a(out_6805),
            .b(out_6811),
            .outp(out_6812)
        );        
        

        logic [WIDTH-1:0] out_6813;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.325)
        ) inst_6813 (
            .outp(out_6813)
        );
        

        logic [WIDTH-1:0] out_6814;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6814 (
            .a(out_14),
            .b(out_6813),
            .outp(out_6814)
        );        
        

        logic [WIDTH-1:0] out_6815;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6815 (
            .a(out_6462),
            .b(out_6814),
            .outp(out_6815)
        );        
        

        logic [WIDTH-1:0] out_6816;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5705)
        ) inst_6816 (
            .outp(out_6816)
        );
        

        logic [WIDTH-1:0] out_6817;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6817 (
            .a(out_3),
            .b(out_6816),
            .outp(out_6817)
        );        
        

        logic [WIDTH-1:0] out_6818;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6818 (
            .a(out_6815),
            .b(out_6817),
            .outp(out_6818)
        );        
        

        logic [WIDTH-1:0] out_6819;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.4705)
        ) inst_6819 (
            .outp(out_6819)
        );
        

        logic [WIDTH-1:0] out_6820;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6820 (
            .a(out_6819),
            .b(out_3),
            .outp(out_6820)
        );        
        

        logic [WIDTH-1:0] out_6821;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6821 (
            .a(out_6818),
            .b(out_6820),
            .outp(out_6821)
        );        
        

        logic [WIDTH-1:0] out_6822;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6822 (
            .a(out_6812),
            .b(out_6821),
            .outp(out_6822)
        );        
        

        logic [WIDTH-1:0] out_6823;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.45)
        ) inst_6823 (
            .outp(out_6823)
        );
        

        logic [WIDTH-1:0] out_6824;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6824 (
            .a(out_14),
            .b(out_6823),
            .outp(out_6824)
        );        
        

        logic [WIDTH-1:0] out_6825;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6825 (
            .a(out_6820),
            .b(out_6824),
            .outp(out_6825)
        );        
        

        logic [WIDTH-1:0] out_6826;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6826 (
            .a(out_6657),
            .b(out_14),
            .outp(out_6826)
        );        
        

        logic [WIDTH-1:0] out_6827;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6827 (
            .a(out_6825),
            .b(out_6826),
            .outp(out_6827)
        );        
        

        logic [WIDTH-1:0] out_6828;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.1205)
        ) inst_6828 (
            .outp(out_6828)
        );
        

        logic [WIDTH-1:0] out_6829;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6829 (
            .a(out_3),
            .b(out_6828),
            .outp(out_6829)
        );        
        

        logic [WIDTH-1:0] out_6830;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6830 (
            .a(out_6827),
            .b(out_6829),
            .outp(out_6830)
        );        
        

        logic [WIDTH-1:0] out_6831;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6831 (
            .in(out_6781),
            .outp(out_6831)
        );
        

        logic [WIDTH-1:0] out_6832;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8955)
        ) inst_6832 (
            .outp(out_6832)
        );
        

        logic [WIDTH-1:0] out_6833;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6833 (
            .a(out_3),
            .b(out_6832),
            .outp(out_6833)
        );        
        

        logic [WIDTH-1:0] out_6834;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6834 (
            .in(out_6833),
            .outp(out_6834)
        );
        

        logic [WIDTH-1:0] out_6835;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6835 (
            .a(out_6831),
            .b(out_6834),
            .outp(out_6835)
        );        
        

        logic [WIDTH-1:0] out_6836;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6836 (
            .in(out_6835),
            .outp(out_6836)
        );
        

        logic [WIDTH-1:0] out_6837;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6837 (
            .a(out_460),
            .b(out_6836),
            .outp(out_6837)
        );        
        

        logic [WIDTH-1:0] out_6838;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6838 (
            .a(out_6836),
            .b(out_9),
            .outp(out_6838)
        );        
        

        logic [WIDTH-1:0] out_6839;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6839 (
            .a(out_6837),
            .b(out_6838),
            .outp(out_6839)
        );        
        

        logic [WIDTH-1:0] out_6840;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.6455)
        ) inst_6840 (
            .outp(out_6840)
        );
        

        logic [WIDTH-1:0] out_6841;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6841 (
            .a(out_3),
            .b(out_6840),
            .outp(out_6841)
        );        
        

        logic [WIDTH-1:0] out_6842;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6842 (
            .in(out_6841),
            .outp(out_6842)
        );
        

        logic [WIDTH-1:0] out_6843;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6843 (
            .a(out_6831),
            .b(out_6842),
            .outp(out_6843)
        );        
        

        logic [WIDTH-1:0] out_6844;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6844 (
            .in(out_6843),
            .outp(out_6844)
        );
        

        logic [WIDTH-1:0] out_6845;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6845 (
            .a(out_460),
            .b(out_6844),
            .outp(out_6845)
        );        
        

        logic [WIDTH-1:0] out_6846;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6846 (
            .a(out_6844),
            .b(out_9),
            .outp(out_6846)
        );        
        

        logic [WIDTH-1:0] out_6847;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6847 (
            .a(out_6845),
            .b(out_6846),
            .outp(out_6847)
        );        
        

        logic [WIDTH-1:0] out_6848;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6848 (
            .a(out_6839),
            .b(out_6847),
            .outp(out_6848)
        );        
        

        logic [WIDTH-1:0] out_6849;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6849 (
            .a(out_6830),
            .b(out_6848),
            .outp(out_6849)
        );        
        

        logic [WIDTH-1:0] out_6850;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6850 (
            .a(out_6822),
            .b(out_6849),
            .outp(out_6850)
        );        
        

        logic [WIDTH-1:0] out_6851;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.6205)
        ) inst_6851 (
            .outp(out_6851)
        );
        

        logic [WIDTH-1:0] out_6852;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6852 (
            .a(out_3),
            .b(out_6851),
            .outp(out_6852)
        );        
        

        logic [WIDTH-1:0] out_6853;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6853 (
            .a(out_6729),
            .b(out_6852),
            .outp(out_6853)
        );        
        

        logic [WIDTH-1:0] out_6854;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5205)
        ) inst_6854 (
            .outp(out_6854)
        );
        

        logic [WIDTH-1:0] out_6855;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6855 (
            .a(out_6854),
            .b(out_3),
            .outp(out_6855)
        );        
        

        logic [WIDTH-1:0] out_6856;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6856 (
            .a(out_6853),
            .b(out_6855),
            .outp(out_6856)
        );        
        

        logic [WIDTH-1:0] out_6857;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6857 (
            .a(out_6850),
            .b(out_6856),
            .outp(out_6857)
        );        
        

        logic [WIDTH-1:0] out_6858;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6858 (
            .a(out_6462),
            .b(out_6477),
            .outp(out_6858)
        );        
        

        logic [WIDTH-1:0] out_6859;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.1705)
        ) inst_6859 (
            .outp(out_6859)
        );
        

        logic [WIDTH-1:0] out_6860;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6860 (
            .a(out_3),
            .b(out_6859),
            .outp(out_6860)
        );        
        

        logic [WIDTH-1:0] out_6861;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6861 (
            .a(out_6858),
            .b(out_6860),
            .outp(out_6861)
        );        
        

        logic [WIDTH-1:0] out_6862;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.0705)
        ) inst_6862 (
            .outp(out_6862)
        );
        

        logic [WIDTH-1:0] out_6863;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6863 (
            .a(out_6862),
            .b(out_3),
            .outp(out_6863)
        );        
        

        logic [WIDTH-1:0] out_6864;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6864 (
            .a(out_6861),
            .b(out_6863),
            .outp(out_6864)
        );        
        

        logic [WIDTH-1:0] out_6865;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6865 (
            .a(out_6857),
            .b(out_6864),
            .outp(out_6865)
        );        
        

        logic [WIDTH-1:0] out_6866;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6866 (
            .a(out_6509),
            .b(out_6852),
            .outp(out_6866)
        );        
        

        logic [WIDTH-1:0] out_6867;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6867 (
            .a(out_6866),
            .b(out_6863),
            .outp(out_6867)
        );        
        

        logic [WIDTH-1:0] out_6868;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6868 (
            .a(out_6867),
            .b(out_6726),
            .outp(out_6868)
        );        
        

        logic [WIDTH-1:0] out_6869;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.3455)
        ) inst_6869 (
            .outp(out_6869)
        );
        

        logic [WIDTH-1:0] out_6870;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6870 (
            .a(out_3),
            .b(out_6869),
            .outp(out_6870)
        );        
        

        logic [WIDTH-1:0] out_6871;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6871 (
            .in(out_6870),
            .outp(out_6871)
        );
        

        logic [WIDTH-1:0] out_6872;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6872 (
            .a(out_6498),
            .b(out_6871),
            .outp(out_6872)
        );        
        

        logic [WIDTH-1:0] out_6873;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6873 (
            .in(out_6872),
            .outp(out_6873)
        );
        

        logic [WIDTH-1:0] out_6874;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6874 (
            .a(out_9),
            .b(out_6873),
            .outp(out_6874)
        );        
        

        logic [WIDTH-1:0] out_6875;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6875 (
            .a(out_6868),
            .b(out_6874),
            .outp(out_6875)
        );        
        

        logic [WIDTH-1:0] out_6876;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6876 (
            .a(out_6873),
            .b(out_21),
            .outp(out_6876)
        );        
        

        logic [WIDTH-1:0] out_6877;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6877 (
            .a(out_6875),
            .b(out_6876),
            .outp(out_6877)
        );        
        

        logic [WIDTH-1:0] out_6878;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6878 (
            .a(out_6865),
            .b(out_6877),
            .outp(out_6878)
        );        
        

        logic [WIDTH-1:0] out_6879;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.825)
        ) inst_6879 (
            .outp(out_6879)
        );
        

        logic [WIDTH-1:0] out_6880;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6880 (
            .a(out_6879),
            .b(out_14),
            .outp(out_6880)
        );        
        

        logic [WIDTH-1:0] out_6881;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.4085)
        ) inst_6881 (
            .outp(out_6881)
        );
        

        logic [WIDTH-1:0] out_6882;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6882 (
            .a(out_3),
            .b(out_6881),
            .outp(out_6882)
        );        
        

        logic [WIDTH-1:0] out_6883;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6883 (
            .a(out_6880),
            .b(out_6882),
            .outp(out_6883)
        );        
        

        logic [WIDTH-1:0] out_6884;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.9085)
        ) inst_6884 (
            .outp(out_6884)
        );
        

        logic [WIDTH-1:0] out_6885;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6885 (
            .a(out_6884),
            .b(out_3),
            .outp(out_6885)
        );        
        

        logic [WIDTH-1:0] out_6886;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6886 (
            .a(out_6883),
            .b(out_6885),
            .outp(out_6886)
        );        
        

        logic [WIDTH-1:0] out_6887;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.915)
        ) inst_6887 (
            .outp(out_6887)
        );
        

        logic [WIDTH-1:0] out_6888;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6888 (
            .a(out_14),
            .b(out_6887),
            .outp(out_6888)
        );        
        

        logic [WIDTH-1:0] out_6889;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6889 (
            .a(out_6886),
            .b(out_6888),
            .outp(out_6889)
        );        
        

        logic [WIDTH-1:0] out_6890;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.51875)
        ) inst_6890 (
            .outp(out_6890)
        );
        

        logic [WIDTH-1:0] out_6891;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6891 (
            .a(out_553),
            .b(out_6890),
            .outp(out_6891)
        );        
        

        logic [WIDTH-1:0] out_6892;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.23609)
        ) inst_6892 (
            .outp(out_6892)
        );
        

        logic [WIDTH-1:0] out_6893;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6893 (
            .a(out_559),
            .b(out_6892),
            .outp(out_6893)
        );        
        

        logic [WIDTH-1:0] out_6894;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6894 (
            .a(out_556),
            .b(out_6893),
            .outp(out_6894)
        );        
        

        logic [WIDTH-1:0] out_6895;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6895 (
            .a(out_6891),
            .b(out_6894),
            .outp(out_6895)
        );        
        

        logic [WIDTH-1:0] out_6896;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.57609)
        ) inst_6896 (
            .outp(out_6896)
        );
        

        logic [WIDTH-1:0] out_6897;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6897 (
            .a(out_6896),
            .b(out_2653),
            .outp(out_6897)
        );        
        

        logic [WIDTH-1:0] out_6898;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6898 (
            .a(out_6895),
            .b(out_6897),
            .outp(out_6898)
        );        
        

        logic [WIDTH-1:0] out_6899;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6899 (
            .a(out_2653),
            .b(out_6896),
            .outp(out_6899)
        );        
        

        logic [WIDTH-1:0] out_6900;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6900 (
            .a(out_6893),
            .b(out_556),
            .outp(out_6900)
        );        
        

        logic [WIDTH-1:0] out_6901;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6901 (
            .a(out_6899),
            .b(out_6900),
            .outp(out_6901)
        );        
        

        logic [WIDTH-1:0] out_6902;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6902 (
            .a(out_6890),
            .b(out_553),
            .outp(out_6902)
        );        
        

        logic [WIDTH-1:0] out_6903;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6903 (
            .a(out_6901),
            .b(out_6902),
            .outp(out_6903)
        );        
        

        logic [WIDTH-1:0] out_6904;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6904 (
            .a(out_6898),
            .b(out_6903),
            .outp(out_6904)
        );        
        

        logic [WIDTH-1:0] out_6905;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6905 (
            .in(out_6904),
            .outp(out_6905)
        );
        

        logic [WIDTH-1:0] out_6906;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.875)
        ) inst_6906 (
            .outp(out_6906)
        );
        

        logic [WIDTH-1:0] out_6907;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6907 (
            .a(out_14),
            .b(out_6906),
            .outp(out_6907)
        );        
        

        logic [WIDTH-1:0] out_6908;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6908 (
            .in(out_6907),
            .outp(out_6908)
        );
        

        logic [WIDTH-1:0] out_6909;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.1335)
        ) inst_6909 (
            .outp(out_6909)
        );
        

        logic [WIDTH-1:0] out_6910;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6910 (
            .a(out_3),
            .b(out_6909),
            .outp(out_6910)
        );        
        

        logic [WIDTH-1:0] out_6911;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6911 (
            .in(out_6910),
            .outp(out_6911)
        );
        

        logic [WIDTH-1:0] out_6912;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6912 (
            .a(out_6908),
            .b(out_6911),
            .outp(out_6912)
        );        
        

        logic [WIDTH-1:0] out_6913;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6913 (
            .in(out_6912),
            .outp(out_6913)
        );
        

        logic [WIDTH-1:0] out_6914;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6914 (
            .a(out_9),
            .b(out_6913),
            .outp(out_6914)
        );        
        

        logic [WIDTH-1:0] out_6915;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6915 (
            .a(out_6905),
            .b(out_6914),
            .outp(out_6915)
        );        
        

        logic [WIDTH-1:0] out_6916;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6916 (
            .a(out_6913),
            .b(out_21),
            .outp(out_6916)
        );        
        

        logic [WIDTH-1:0] out_6917;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6917 (
            .a(out_6915),
            .b(out_6916),
            .outp(out_6917)
        );        
        

        logic [WIDTH-1:0] out_6918;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6918 (
            .a(out_6889),
            .b(out_6917),
            .outp(out_6918)
        );        
        

        logic [WIDTH-1:0] out_6919;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6919 (
            .a(out_6918),
            .b(out_6916),
            .outp(out_6919)
        );        
        

        logic [WIDTH-1:0] out_6920;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6920 (
            .a(out_6878),
            .b(out_6919),
            .outp(out_6920)
        );        
        

        logic [WIDTH-1:0] out_6921;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.95)
        ) inst_6921 (
            .outp(out_6921)
        );
        

        logic [WIDTH-1:0] out_6922;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6922 (
            .a(out_14),
            .b(out_6921),
            .outp(out_6922)
        );        
        

        logic [WIDTH-1:0] out_6923;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.6)
        ) inst_6923 (
            .outp(out_6923)
        );
        

        logic [WIDTH-1:0] out_6924;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6924 (
            .a(out_6923),
            .b(out_14),
            .outp(out_6924)
        );        
        

        logic [WIDTH-1:0] out_6925;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6925 (
            .a(out_6922),
            .b(out_6924),
            .outp(out_6925)
        );        
        

        logic [WIDTH-1:0] out_6926;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.7585)
        ) inst_6926 (
            .outp(out_6926)
        );
        

        logic [WIDTH-1:0] out_6927;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6927 (
            .a(out_3),
            .b(out_6926),
            .outp(out_6927)
        );        
        

        logic [WIDTH-1:0] out_6928;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6928 (
            .a(out_6925),
            .b(out_6927),
            .outp(out_6928)
        );        
        

        logic [WIDTH-1:0] out_6929;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.6585)
        ) inst_6929 (
            .outp(out_6929)
        );
        

        logic [WIDTH-1:0] out_6930;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6930 (
            .a(out_6929),
            .b(out_3),
            .outp(out_6930)
        );        
        

        logic [WIDTH-1:0] out_6931;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6931 (
            .a(out_6928),
            .b(out_6930),
            .outp(out_6931)
        );        
        

        logic [WIDTH-1:0] out_6932;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6932 (
            .a(out_6920),
            .b(out_6931),
            .outp(out_6932)
        );        
        

        logic [WIDTH-1:0] out_6933;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.5085)
        ) inst_6933 (
            .outp(out_6933)
        );
        

        logic [WIDTH-1:0] out_6934;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6934 (
            .a(out_3),
            .b(out_6933),
            .outp(out_6934)
        );        
        

        logic [WIDTH-1:0] out_6935;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6935 (
            .a(out_6925),
            .b(out_6934),
            .outp(out_6935)
        );        
        

        logic [WIDTH-1:0] out_6936;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.4085)
        ) inst_6936 (
            .outp(out_6936)
        );
        

        logic [WIDTH-1:0] out_6937;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6937 (
            .a(out_6936),
            .b(out_3),
            .outp(out_6937)
        );        
        

        logic [WIDTH-1:0] out_6938;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6938 (
            .a(out_6935),
            .b(out_6937),
            .outp(out_6938)
        );        
        

        logic [WIDTH-1:0] out_6939;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6939 (
            .a(out_6932),
            .b(out_6938),
            .outp(out_6939)
        );        
        

        logic [WIDTH-1:0] out_6940;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.125)
        ) inst_6940 (
            .outp(out_6940)
        );
        

        logic [WIDTH-1:0] out_6941;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6941 (
            .a(out_14),
            .b(out_6940),
            .outp(out_6941)
        );        
        

        logic [WIDTH-1:0] out_6942;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6942 (
            .a(out_6924),
            .b(out_6941),
            .outp(out_6942)
        );        
        

        logic [WIDTH-1:0] out_6943;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.2585)
        ) inst_6943 (
            .outp(out_6943)
        );
        

        logic [WIDTH-1:0] out_6944;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6944 (
            .a(out_3),
            .b(out_6943),
            .outp(out_6944)
        );        
        

        logic [WIDTH-1:0] out_6945;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6945 (
            .a(out_6942),
            .b(out_6944),
            .outp(out_6945)
        );        
        

        logic [WIDTH-1:0] out_6946;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.1585)
        ) inst_6946 (
            .outp(out_6946)
        );
        

        logic [WIDTH-1:0] out_6947;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6947 (
            .a(out_6946),
            .b(out_3),
            .outp(out_6947)
        );        
        

        logic [WIDTH-1:0] out_6948;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6948 (
            .a(out_6945),
            .b(out_6947),
            .outp(out_6948)
        );        
        

        logic [WIDTH-1:0] out_6949;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6949 (
            .a(out_6939),
            .b(out_6948),
            .outp(out_6949)
        );        
        

        logic [WIDTH-1:0] out_6950;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.25)
        ) inst_6950 (
            .outp(out_6950)
        );
        

        logic [WIDTH-1:0] out_6951;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6951 (
            .a(out_14),
            .b(out_6950),
            .outp(out_6951)
        );        
        

        logic [WIDTH-1:0] out_6952;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6952 (
            .a(out_6947),
            .b(out_6951),
            .outp(out_6952)
        );        
        

        logic [WIDTH-1:0] out_6953;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.95)
        ) inst_6953 (
            .outp(out_6953)
        );
        

        logic [WIDTH-1:0] out_6954;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6954 (
            .a(out_6953),
            .b(out_14),
            .outp(out_6954)
        );        
        

        logic [WIDTH-1:0] out_6955;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6955 (
            .a(out_6952),
            .b(out_6954),
            .outp(out_6955)
        );        
        

        logic [WIDTH-1:0] out_6956;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.8085)
        ) inst_6956 (
            .outp(out_6956)
        );
        

        logic [WIDTH-1:0] out_6957;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6957 (
            .a(out_3),
            .b(out_6956),
            .outp(out_6957)
        );        
        

        logic [WIDTH-1:0] out_6958;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6958 (
            .a(out_6955),
            .b(out_6957),
            .outp(out_6958)
        );        
        

        logic [WIDTH-1:0] out_6959;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6959 (
            .in(out_6922),
            .outp(out_6959)
        );
        

        logic [WIDTH-1:0] out_6960;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.5835)
        ) inst_6960 (
            .outp(out_6960)
        );
        

        logic [WIDTH-1:0] out_6961;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6961 (
            .a(out_3),
            .b(out_6960),
            .outp(out_6961)
        );        
        

        logic [WIDTH-1:0] out_6962;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6962 (
            .in(out_6961),
            .outp(out_6962)
        );
        

        logic [WIDTH-1:0] out_6963;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6963 (
            .a(out_6959),
            .b(out_6962),
            .outp(out_6963)
        );        
        

        logic [WIDTH-1:0] out_6964;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6964 (
            .in(out_6963),
            .outp(out_6964)
        );
        

        logic [WIDTH-1:0] out_6965;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6965 (
            .a(out_460),
            .b(out_6964),
            .outp(out_6965)
        );        
        

        logic [WIDTH-1:0] out_6966;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6966 (
            .a(out_6964),
            .b(out_9),
            .outp(out_6966)
        );        
        

        logic [WIDTH-1:0] out_6967;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6967 (
            .a(out_6965),
            .b(out_6966),
            .outp(out_6967)
        );        
        

        logic [WIDTH-1:0] out_6968;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.3335)
        ) inst_6968 (
            .outp(out_6968)
        );
        

        logic [WIDTH-1:0] out_6969;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6969 (
            .a(out_3),
            .b(out_6968),
            .outp(out_6969)
        );        
        

        logic [WIDTH-1:0] out_6970;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6970 (
            .in(out_6969),
            .outp(out_6970)
        );
        

        logic [WIDTH-1:0] out_6971;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6971 (
            .a(out_6959),
            .b(out_6970),
            .outp(out_6971)
        );        
        

        logic [WIDTH-1:0] out_6972;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6972 (
            .in(out_6971),
            .outp(out_6972)
        );
        

        logic [WIDTH-1:0] out_6973;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6973 (
            .a(out_460),
            .b(out_6972),
            .outp(out_6973)
        );        
        

        logic [WIDTH-1:0] out_6974;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6974 (
            .a(out_6972),
            .b(out_9),
            .outp(out_6974)
        );        
        

        logic [WIDTH-1:0] out_6975;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6975 (
            .a(out_6973),
            .b(out_6974),
            .outp(out_6975)
        );        
        

        logic [WIDTH-1:0] out_6976;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6976 (
            .a(out_6967),
            .b(out_6975),
            .outp(out_6976)
        );        
        

        logic [WIDTH-1:0] out_6977;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6977 (
            .a(out_6958),
            .b(out_6976),
            .outp(out_6977)
        );        
        

        logic [WIDTH-1:0] out_6978;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6978 (
            .a(out_6949),
            .b(out_6977),
            .outp(out_6978)
        );        
        

        logic [WIDTH-1:0] out_6979;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6979 (
            .a(out_4460),
            .b(out_5137),
            .outp(out_6979)
        );        
        

        logic [WIDTH-1:0] out_6980;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6980 (
            .in(out_5142),
            .outp(out_6980)
        );
        

        logic [WIDTH-1:0] out_6981;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6981 (
            .a(out_6979),
            .b(out_6980),
            .outp(out_6981)
        );        
        

        logic [WIDTH-1:0] out_6982;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6982 (
            .a(out_6978),
            .b(out_6981),
            .outp(out_6982)
        );        
        

        logic [WIDTH-1:0] out_6983;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6983 (
            .a(out_4464),
            .b(out_6980),
            .outp(out_6983)
        );        
        

        logic [WIDTH-1:0] out_6984;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.466)
        ) inst_6984 (
            .outp(out_6984)
        );
        

        logic [WIDTH-1:0] out_6985;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6985 (
            .a(out_131),
            .b(out_6984),
            .outp(out_6985)
        );        
        

        logic [WIDTH-1:0] out_6986;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6986 (
            .a(out_6985),
            .b(out_127),
            .outp(out_6986)
        );        
        

        logic [WIDTH-1:0] out_6987;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6987 (
            .a(out_6983),
            .b(out_6986),
            .outp(out_6987)
        );        
        

        logic [WIDTH-1:0] out_6988;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6988 (
            .a(out_6982),
            .b(out_6987),
            .outp(out_6988)
        );        
        

        logic [WIDTH-1:0] out_6989;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6989 (
            .a(out_4473),
            .b(out_5142),
            .outp(out_6989)
        );        
        

        logic [WIDTH-1:0] out_6990;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6990 (
            .in(out_6986),
            .outp(out_6990)
        );
        

        logic [WIDTH-1:0] out_6991;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6991 (
            .a(out_6989),
            .b(out_6990),
            .outp(out_6991)
        );        
        

        logic [WIDTH-1:0] out_6992;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6992 (
            .a(out_6988),
            .b(out_6991),
            .outp(out_6992)
        );        
        

        logic [WIDTH-1:0] out_6993;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.09)
        ) inst_6993 (
            .outp(out_6993)
        );
        

        logic [WIDTH-1:0] out_6994;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6994 (
            .a(out_6993),
            .b(out_3),
            .outp(out_6994)
        );        
        

        logic [WIDTH-1:0] out_6995;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6995 (
            .a(out_4931),
            .b(out_6994),
            .outp(out_6995)
        );        
        

        logic [WIDTH-1:0] out_6996;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.19)
        ) inst_6996 (
            .outp(out_6996)
        );
        

        logic [WIDTH-1:0] out_6997;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6997 (
            .a(out_6996),
            .b(out_3),
            .outp(out_6997)
        );        
        

        logic [WIDTH-1:0] out_6998;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6998 (
            .in(out_6997),
            .outp(out_6998)
        );
        

        logic [WIDTH-1:0] out_6999;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_6999 (
            .a(out_6995),
            .b(out_6998),
            .outp(out_6999)
        );        
        

        logic [WIDTH-1:0] out_7000;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7000 (
            .a(out_6992),
            .b(out_6999),
            .outp(out_7000)
        );        
        

        logic [WIDTH-1:0] out_7001;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.16429)
        ) inst_7001 (
            .outp(out_7001)
        );
        

        logic [WIDTH-1:0] out_7002;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7002 (
            .a(out_7001),
            .b(out_3),
            .outp(out_7002)
        );        
        

        logic [WIDTH-1:0] out_7003;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7003 (
            .a(out_7002),
            .b(out_1495),
            .outp(out_7003)
        );        
        

        logic [WIDTH-1:0] out_7004;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7004 (
            .in(out_7003),
            .outp(out_7004)
        );
        

        logic [WIDTH-1:0] out_7005;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7005 (
            .a(out_4420),
            .b(out_7004),
            .outp(out_7005)
        );        
        

        logic [WIDTH-1:0] out_7006;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7006 (
            .in(out_7005),
            .outp(out_7006)
        );
        

        logic [WIDTH-1:0] out_7007;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7007 (
            .a(out_9),
            .b(out_7006),
            .outp(out_7007)
        );        
        

        logic [WIDTH-1:0] out_7008;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7008 (
            .a(out_7006),
            .b(out_21),
            .outp(out_7008)
        );        
        

        logic [WIDTH-1:0] out_7009;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7009 (
            .a(out_7007),
            .b(out_7008),
            .outp(out_7009)
        );        
        

        logic [WIDTH-1:0] out_7010;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7010 (
            .a(out_7000),
            .b(out_7009),
            .outp(out_7010)
        );        
        

        logic [WIDTH-1:0] out_7011;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7011 (
            .a(out_4409),
            .b(out_4542),
            .outp(out_7011)
        );        
        

        logic [WIDTH-1:0] out_7012;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7012 (
            .in(out_5346),
            .outp(out_7012)
        );
        

        logic [WIDTH-1:0] out_7013;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7013 (
            .a(out_7011),
            .b(out_7012),
            .outp(out_7013)
        );        
        

        logic [WIDTH-1:0] out_7014;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7014 (
            .a(out_4565),
            .b(out_4420),
            .outp(out_7014)
        );        
        

        logic [WIDTH-1:0] out_7015;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7015 (
            .in(out_7014),
            .outp(out_7015)
        );
        

        logic [WIDTH-1:0] out_7016;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7016 (
            .a(out_7015),
            .b(out_21),
            .outp(out_7016)
        );        
        

        logic [WIDTH-1:0] out_7017;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.2175)
        ) inst_7017 (
            .outp(out_7017)
        );
        

        logic [WIDTH-1:0] out_7018;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7018 (
            .a(out_7017),
            .b(out_556),
            .outp(out_7018)
        );        
        

        logic [WIDTH-1:0] out_7019;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7019 (
            .a(out_7018),
            .b(out_559),
            .outp(out_7019)
        );        
        

        logic [WIDTH-1:0] out_7020;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7020 (
            .a(out_4425),
            .b(out_7019),
            .outp(out_7020)
        );        
        

        logic [WIDTH-1:0] out_7021;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5925)
        ) inst_7021 (
            .outp(out_7021)
        );
        

        logic [WIDTH-1:0] out_7022;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7022 (
            .a(out_7021),
            .b(out_556),
            .outp(out_7022)
        );        
        

        logic [WIDTH-1:0] out_7023;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7023 (
            .a(out_7022),
            .b(out_566),
            .outp(out_7023)
        );        
        

        logic [WIDTH-1:0] out_7024;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7024 (
            .in(out_7023),
            .outp(out_7024)
        );
        

        logic [WIDTH-1:0] out_7025;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7025 (
            .a(out_7020),
            .b(out_7024),
            .outp(out_7025)
        );        
        

        logic [WIDTH-1:0] out_7026;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5925)
        ) inst_7026 (
            .outp(out_7026)
        );
        

        logic [WIDTH-1:0] out_7027;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7027 (
            .a(out_7026),
            .b(out_556),
            .outp(out_7027)
        );        
        

        logic [WIDTH-1:0] out_7028;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7028 (
            .a(out_7027),
            .b(out_566),
            .outp(out_7028)
        );        
        

        logic [WIDTH-1:0] out_7029;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7029 (
            .a(out_4436),
            .b(out_7028),
            .outp(out_7029)
        );        
        

        logic [WIDTH-1:0] out_7030;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7030 (
            .a(out_559),
            .b(out_7018),
            .outp(out_7030)
        );        
        

        logic [WIDTH-1:0] out_7031;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7031 (
            .a(out_7029),
            .b(out_7030),
            .outp(out_7031)
        );        
        

        logic [WIDTH-1:0] out_7032;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7032 (
            .a(out_7025),
            .b(out_7031),
            .outp(out_7032)
        );        
        

        logic [WIDTH-1:0] out_7033;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7033 (
            .in(out_7032),
            .outp(out_7033)
        );
        

        logic [WIDTH-1:0] out_7034;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7034 (
            .a(out_7016),
            .b(out_7033),
            .outp(out_7034)
        );        
        

        logic [WIDTH-1:0] out_7035;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7035 (
            .a(out_9),
            .b(out_7015),
            .outp(out_7035)
        );        
        

        logic [WIDTH-1:0] out_7036;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7036 (
            .a(out_7034),
            .b(out_7035),
            .outp(out_7036)
        );        
        

        logic [WIDTH-1:0] out_7037;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7037 (
            .a(out_7013),
            .b(out_7036),
            .outp(out_7037)
        );        
        

        logic [WIDTH-1:0] out_7038;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7038 (
            .a(out_7016),
            .b(out_7037),
            .outp(out_7038)
        );        
        

        logic [WIDTH-1:0] out_7039;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7039 (
            .a(out_7010),
            .b(out_7038),
            .outp(out_7039)
        );        
        

        logic [WIDTH-1:0] out_7040;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7040 (
            .a(out_2782),
            .b(out_4580),
            .outp(out_7040)
        );        
        

        logic [WIDTH-1:0] out_7041;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7041 (
            .a(out_7040),
            .b(out_4419),
            .outp(out_7041)
        );        
        

        logic [WIDTH-1:0] out_7042;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.55)
        ) inst_7042 (
            .outp(out_7042)
        );
        

        logic [WIDTH-1:0] out_7043;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7043 (
            .a(out_7042),
            .b(out_3),
            .outp(out_7043)
        );        
        

        logic [WIDTH-1:0] out_7044;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7044 (
            .in(out_7043),
            .outp(out_7044)
        );
        

        logic [WIDTH-1:0] out_7045;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7045 (
            .a(out_7041),
            .b(out_7044),
            .outp(out_7045)
        );        
        

        logic [WIDTH-1:0] out_7046;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7046 (
            .a(out_7039),
            .b(out_7045),
            .outp(out_7046)
        );        
        

        logic [WIDTH-1:0] out_7047;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(7.9)
        ) inst_7047 (
            .outp(out_7047)
        );
        

        logic [WIDTH-1:0] out_7048;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7048 (
            .a(out_7047),
            .b(out_3),
            .outp(out_7048)
        );        
        

        logic [WIDTH-1:0] out_7049;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7049 (
            .a(out_4775),
            .b(out_7048),
            .outp(out_7049)
        );        
        

        logic [WIDTH-1:0] out_7050;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(8.0)
        ) inst_7050 (
            .outp(out_7050)
        );
        

        logic [WIDTH-1:0] out_7051;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7051 (
            .a(out_7050),
            .b(out_3),
            .outp(out_7051)
        );        
        

        logic [WIDTH-1:0] out_7052;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7052 (
            .in(out_7051),
            .outp(out_7052)
        );
        

        logic [WIDTH-1:0] out_7053;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7053 (
            .a(out_7049),
            .b(out_7052),
            .outp(out_7053)
        );        
        

        logic [WIDTH-1:0] out_7054;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7054 (
            .a(out_7046),
            .b(out_7053),
            .outp(out_7054)
        );        
        

        logic [WIDTH-1:0] out_7055;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7055 (
            .a(out_2782),
            .b(out_4590),
            .outp(out_7055)
        );        
        

        logic [WIDTH-1:0] out_7056;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7056 (
            .a(out_7055),
            .b(out_4641),
            .outp(out_7056)
        );        
        

        logic [WIDTH-1:0] out_7057;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7057 (
            .a(out_7056),
            .b(out_7052),
            .outp(out_7057)
        );        
        

        logic [WIDTH-1:0] out_7058;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7058 (
            .a(out_2790),
            .b(out_4420),
            .outp(out_7058)
        );        
        

        logic [WIDTH-1:0] out_7059;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7059 (
            .in(out_7058),
            .outp(out_7059)
        );
        

        logic [WIDTH-1:0] out_7060;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7060 (
            .a(out_9),
            .b(out_7059),
            .outp(out_7060)
        );        
        

        logic [WIDTH-1:0] out_7061;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7061 (
            .a(out_7057),
            .b(out_7060),
            .outp(out_7061)
        );        
        

        logic [WIDTH-1:0] out_7062;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7062 (
            .a(out_7059),
            .b(out_21),
            .outp(out_7062)
        );        
        

        logic [WIDTH-1:0] out_7063;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7063 (
            .a(out_7061),
            .b(out_7062),
            .outp(out_7063)
        );        
        

        logic [WIDTH-1:0] out_7064;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7064 (
            .a(out_7054),
            .b(out_7063),
            .outp(out_7064)
        );        
        

        logic [WIDTH-1:0] out_7065;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7065 (
            .a(out_6924),
            .b(out_6448),
            .outp(out_7065)
        );        
        

        logic [WIDTH-1:0] out_7066;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.121)
        ) inst_7066 (
            .outp(out_7066)
        );
        

        logic [WIDTH-1:0] out_7067;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7067 (
            .a(out_7066),
            .b(out_3),
            .outp(out_7067)
        );        
        

        logic [WIDTH-1:0] out_7068;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7068 (
            .a(out_7065),
            .b(out_7067),
            .outp(out_7068)
        );        
        

        logic [WIDTH-1:0] out_7069;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.846)
        ) inst_7069 (
            .outp(out_7069)
        );
        

        logic [WIDTH-1:0] out_7070;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7070 (
            .a(out_3),
            .b(out_7069),
            .outp(out_7070)
        );        
        

        logic [WIDTH-1:0] out_7071;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7071 (
            .a(out_7068),
            .b(out_7070),
            .outp(out_7071)
        );        
        

        logic [WIDTH-1:0] out_7072;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.846)
        ) inst_7072 (
            .outp(out_7072)
        );
        

        logic [WIDTH-1:0] out_7073;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7073 (
            .a(out_7072),
            .b(out_3),
            .outp(out_7073)
        );        
        

        logic [WIDTH-1:0] out_7074;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7074 (
            .in(out_7073),
            .outp(out_7074)
        );
        

        logic [WIDTH-1:0] out_7075;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7075 (
            .a(out_6908),
            .b(out_7074),
            .outp(out_7075)
        );        
        

        logic [WIDTH-1:0] out_7076;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7076 (
            .in(out_7075),
            .outp(out_7076)
        );
        

        logic [WIDTH-1:0] out_7077;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7077 (
            .a(out_9),
            .b(out_7076),
            .outp(out_7077)
        );        
        

        logic [WIDTH-1:0] out_7078;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7078 (
            .a(out_7071),
            .b(out_7077),
            .outp(out_7078)
        );        
        

        logic [WIDTH-1:0] out_7079;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7079 (
            .a(out_7076),
            .b(out_21),
            .outp(out_7079)
        );        
        

        logic [WIDTH-1:0] out_7080;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7080 (
            .a(out_7078),
            .b(out_7079),
            .outp(out_7080)
        );        
        

        logic [WIDTH-1:0] out_7081;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7081 (
            .a(out_7064),
            .b(out_7080),
            .outp(out_7081)
        );        
        

        logic [WIDTH-1:0] out_7082;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7082 (
            .a(out_6880),
            .b(out_6888),
            .outp(out_7082)
        );        
        

        logic [WIDTH-1:0] out_7083;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.496)
        ) inst_7083 (
            .outp(out_7083)
        );
        

        logic [WIDTH-1:0] out_7084;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7084 (
            .a(out_3),
            .b(out_7083),
            .outp(out_7084)
        );        
        

        logic [WIDTH-1:0] out_7085;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7085 (
            .a(out_7082),
            .b(out_7084),
            .outp(out_7085)
        );        
        

        logic [WIDTH-1:0] out_7086;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.996)
        ) inst_7086 (
            .outp(out_7086)
        );
        

        logic [WIDTH-1:0] out_7087;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7087 (
            .a(out_7086),
            .b(out_3),
            .outp(out_7087)
        );        
        

        logic [WIDTH-1:0] out_7088;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7088 (
            .a(out_7085),
            .b(out_7087),
            .outp(out_7088)
        );        
        

        logic [WIDTH-1:0] out_7089;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.221)
        ) inst_7089 (
            .outp(out_7089)
        );
        

        logic [WIDTH-1:0] out_7090;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7090 (
            .a(out_3),
            .b(out_7089),
            .outp(out_7090)
        );        
        

        logic [WIDTH-1:0] out_7091;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7091 (
            .in(out_7090),
            .outp(out_7091)
        );
        

        logic [WIDTH-1:0] out_7092;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7092 (
            .a(out_6908),
            .b(out_7091),
            .outp(out_7092)
        );        
        

        logic [WIDTH-1:0] out_7093;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7093 (
            .in(out_7092),
            .outp(out_7093)
        );
        

        logic [WIDTH-1:0] out_7094;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7094 (
            .a(out_7093),
            .b(out_21),
            .outp(out_7094)
        );        
        

        logic [WIDTH-1:0] out_7095;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.16015)
        ) inst_7095 (
            .outp(out_7095)
        );
        

        logic [WIDTH-1:0] out_7096;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7096 (
            .a(out_7095),
            .b(out_559),
            .outp(out_7096)
        );        
        

        logic [WIDTH-1:0] out_7097;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7097 (
            .a(out_556),
            .b(out_7096),
            .outp(out_7097)
        );        
        

        logic [WIDTH-1:0] out_7098;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7098 (
            .a(out_6891),
            .b(out_7097),
            .outp(out_7098)
        );        
        

        logic [WIDTH-1:0] out_7099;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.50015)
        ) inst_7099 (
            .outp(out_7099)
        );
        

        logic [WIDTH-1:0] out_7100;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7100 (
            .a(out_7099),
            .b(out_2653),
            .outp(out_7100)
        );        
        

        logic [WIDTH-1:0] out_7101;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7101 (
            .a(out_7098),
            .b(out_7100),
            .outp(out_7101)
        );        
        

        logic [WIDTH-1:0] out_7102;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7102 (
            .a(out_2653),
            .b(out_7099),
            .outp(out_7102)
        );        
        

        logic [WIDTH-1:0] out_7103;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7103 (
            .a(out_6902),
            .b(out_7102),
            .outp(out_7103)
        );        
        

        logic [WIDTH-1:0] out_7104;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7104 (
            .a(out_7096),
            .b(out_556),
            .outp(out_7104)
        );        
        

        logic [WIDTH-1:0] out_7105;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7105 (
            .a(out_7103),
            .b(out_7104),
            .outp(out_7105)
        );        
        

        logic [WIDTH-1:0] out_7106;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7106 (
            .a(out_7101),
            .b(out_7105),
            .outp(out_7106)
        );        
        

        logic [WIDTH-1:0] out_7107;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7107 (
            .in(out_7106),
            .outp(out_7107)
        );
        

        logic [WIDTH-1:0] out_7108;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7108 (
            .a(out_7094),
            .b(out_7107),
            .outp(out_7108)
        );        
        

        logic [WIDTH-1:0] out_7109;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7109 (
            .a(out_9),
            .b(out_7093),
            .outp(out_7109)
        );        
        

        logic [WIDTH-1:0] out_7110;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7110 (
            .a(out_7108),
            .b(out_7109),
            .outp(out_7110)
        );        
        

        logic [WIDTH-1:0] out_7111;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7111 (
            .a(out_7088),
            .b(out_7110),
            .outp(out_7111)
        );        
        

        logic [WIDTH-1:0] out_7112;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7112 (
            .a(out_7094),
            .b(out_7111),
            .outp(out_7112)
        );        
        

        logic [WIDTH-1:0] out_7113;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7113 (
            .a(out_7081),
            .b(out_7112),
            .outp(out_7113)
        );        
        

        logic [WIDTH-1:0] out_7114;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.588)
        ) inst_7114 (
            .outp(out_7114)
        );
        

        logic [WIDTH-1:0] out_7115;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7115 (
            .a(out_3),
            .b(out_7114),
            .outp(out_7115)
        );        
        

        logic [WIDTH-1:0] out_7116;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7116 (
            .a(out_6924),
            .b(out_7115),
            .outp(out_7116)
        );        
        

        logic [WIDTH-1:0] out_7117;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.488)
        ) inst_7117 (
            .outp(out_7117)
        );
        

        logic [WIDTH-1:0] out_7118;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7118 (
            .a(out_7117),
            .b(out_3),
            .outp(out_7118)
        );        
        

        logic [WIDTH-1:0] out_7119;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7119 (
            .a(out_7116),
            .b(out_7118),
            .outp(out_7119)
        );        
        

        logic [WIDTH-1:0] out_7120;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.15)
        ) inst_7120 (
            .outp(out_7120)
        );
        

        logic [WIDTH-1:0] out_7121;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7121 (
            .a(out_14),
            .b(out_7120),
            .outp(out_7121)
        );        
        

        logic [WIDTH-1:0] out_7122;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7122 (
            .a(out_7119),
            .b(out_7121),
            .outp(out_7122)
        );        
        

        logic [WIDTH-1:0] out_7123;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7123 (
            .a(out_7113),
            .b(out_7122),
            .outp(out_7123)
        );        
        

        logic [WIDTH-1:0] out_7124;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.67571)
        ) inst_7124 (
            .outp(out_7124)
        );
        

        logic [WIDTH-1:0] out_7125;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7125 (
            .a(out_194),
            .b(out_7124),
            .outp(out_7125)
        );        
        

        logic [WIDTH-1:0] out_7126;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7126 (
            .a(out_6924),
            .b(out_7125),
            .outp(out_7126)
        );        
        

        logic [WIDTH-1:0] out_7127;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.12571)
        ) inst_7127 (
            .outp(out_7127)
        );
        

        logic [WIDTH-1:0] out_7128;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7128 (
            .a(out_7127),
            .b(out_194),
            .outp(out_7128)
        );        
        

        logic [WIDTH-1:0] out_7129;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7129 (
            .a(out_7126),
            .b(out_7128),
            .outp(out_7129)
        );        
        

        logic [WIDTH-1:0] out_7130;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7130 (
            .a(out_14),
            .b(out_6923),
            .outp(out_7130)
        );        
        

        logic [WIDTH-1:0] out_7131;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7131 (
            .in(out_7130),
            .outp(out_7131)
        );
        

        logic [WIDTH-1:0] out_7132;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.34464)
        ) inst_7132 (
            .outp(out_7132)
        );
        

        logic [WIDTH-1:0] out_7133;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7133 (
            .a(out_204),
            .b(out_7132),
            .outp(out_7133)
        );        
        

        logic [WIDTH-1:0] out_7134;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7134 (
            .in(out_7133),
            .outp(out_7134)
        );
        

        logic [WIDTH-1:0] out_7135;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7135 (
            .a(out_7131),
            .b(out_7134),
            .outp(out_7135)
        );        
        

        logic [WIDTH-1:0] out_7136;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7136 (
            .in(out_7135),
            .outp(out_7136)
        );
        

        logic [WIDTH-1:0] out_7137;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7137 (
            .a(out_200),
            .b(out_7136),
            .outp(out_7137)
        );        
        

        logic [WIDTH-1:0] out_7138;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7138 (
            .a(out_7129),
            .b(out_7137),
            .outp(out_7138)
        );        
        

        logic [WIDTH-1:0] out_7139;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7139 (
            .in(out_7125),
            .outp(out_7139)
        );
        

        logic [WIDTH-1:0] out_7140;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7140 (
            .a(out_7131),
            .b(out_7139),
            .outp(out_7140)
        );        
        

        logic [WIDTH-1:0] out_7141;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7141 (
            .in(out_7140),
            .outp(out_7141)
        );
        

        logic [WIDTH-1:0] out_7142;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7142 (
            .a(out_7141),
            .b(out_214),
            .outp(out_7142)
        );        
        

        logic [WIDTH-1:0] out_7143;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7143 (
            .a(out_7138),
            .b(out_7142),
            .outp(out_7143)
        );        
        

        logic [WIDTH-1:0] out_7144;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7144 (
            .a(out_7143),
            .b(out_7121),
            .outp(out_7144)
        );        
        

        logic [WIDTH-1:0] out_7145;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7145 (
            .a(out_7123),
            .b(out_7144),
            .outp(out_7145)
        );        
        

        logic [WIDTH-1:0] out_7146;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.363)
        ) inst_7146 (
            .outp(out_7146)
        );
        

        logic [WIDTH-1:0] out_7147;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7147 (
            .a(out_3),
            .b(out_7146),
            .outp(out_7147)
        );        
        

        logic [WIDTH-1:0] out_7148;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7148 (
            .a(out_6924),
            .b(out_7147),
            .outp(out_7148)
        );        
        

        logic [WIDTH-1:0] out_7149;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.263)
        ) inst_7149 (
            .outp(out_7149)
        );
        

        logic [WIDTH-1:0] out_7150;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7150 (
            .a(out_7149),
            .b(out_3),
            .outp(out_7150)
        );        
        

        logic [WIDTH-1:0] out_7151;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7151 (
            .a(out_7148),
            .b(out_7150),
            .outp(out_7151)
        );        
        

        logic [WIDTH-1:0] out_7152;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7152 (
            .a(out_7151),
            .b(out_7121),
            .outp(out_7152)
        );        
        

        logic [WIDTH-1:0] out_7153;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7153 (
            .a(out_7145),
            .b(out_7152),
            .outp(out_7153)
        );        
        

        logic [WIDTH-1:0] out_7154;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.3)
        ) inst_7154 (
            .outp(out_7154)
        );
        

        logic [WIDTH-1:0] out_7155;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7155 (
            .a(out_14),
            .b(out_7154),
            .outp(out_7155)
        );        
        

        logic [WIDTH-1:0] out_7156;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7156 (
            .in(out_7155),
            .outp(out_7156)
        );
        

        logic [WIDTH-1:0] out_7157;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.313)
        ) inst_7157 (
            .outp(out_7157)
        );
        

        logic [WIDTH-1:0] out_7158;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7158 (
            .a(out_3),
            .b(out_7157),
            .outp(out_7158)
        );        
        

        logic [WIDTH-1:0] out_7159;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7159 (
            .in(out_7158),
            .outp(out_7159)
        );
        

        logic [WIDTH-1:0] out_7160;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7160 (
            .a(out_7156),
            .b(out_7159),
            .outp(out_7160)
        );        
        

        logic [WIDTH-1:0] out_7161;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7161 (
            .in(out_7160),
            .outp(out_7161)
        );
        

        logic [WIDTH-1:0] out_7162;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7162 (
            .a(out_7161),
            .b(out_460),
            .outp(out_7162)
        );        
        

        logic [WIDTH-1:0] out_7163;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7163 (
            .a(out_7153),
            .b(out_7162),
            .outp(out_7163)
        );        
        

        logic [WIDTH-1:0] out_7164;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.138)
        ) inst_7164 (
            .outp(out_7164)
        );
        

        logic [WIDTH-1:0] out_7165;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7165 (
            .a(out_3),
            .b(out_7164),
            .outp(out_7165)
        );        
        

        logic [WIDTH-1:0] out_7166;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7166 (
            .a(out_6924),
            .b(out_7165),
            .outp(out_7166)
        );        
        

        logic [WIDTH-1:0] out_7167;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.038)
        ) inst_7167 (
            .outp(out_7167)
        );
        

        logic [WIDTH-1:0] out_7168;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7168 (
            .a(out_7167),
            .b(out_3),
            .outp(out_7168)
        );        
        

        logic [WIDTH-1:0] out_7169;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7169 (
            .a(out_7166),
            .b(out_7168),
            .outp(out_7169)
        );        
        

        logic [WIDTH-1:0] out_7170;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7170 (
            .a(out_7169),
            .b(out_7121),
            .outp(out_7170)
        );        
        

        logic [WIDTH-1:0] out_7171;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7171 (
            .a(out_7163),
            .b(out_7170),
            .outp(out_7171)
        );        
        

        logic [WIDTH-1:0] out_7172;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.7835)
        ) inst_7172 (
            .outp(out_7172)
        );
        

        logic [WIDTH-1:0] out_7173;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7173 (
            .a(out_3),
            .b(out_7172),
            .outp(out_7173)
        );        
        

        logic [WIDTH-1:0] out_7174;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7174 (
            .in(out_7173),
            .outp(out_7174)
        );
        

        logic [WIDTH-1:0] out_7175;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7175 (
            .a(out_7174),
            .b(out_6908),
            .outp(out_7175)
        );        
        

        logic [WIDTH-1:0] out_7176;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7176 (
            .in(out_7175),
            .outp(out_7176)
        );
        

        logic [WIDTH-1:0] out_7177;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7177 (
            .a(out_7176),
            .b(out_21),
            .outp(out_7177)
        );        
        

        logic [WIDTH-1:0] out_7178;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7178 (
            .a(out_9),
            .b(out_7176),
            .outp(out_7178)
        );        
        

        logic [WIDTH-1:0] out_7179;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7179 (
            .a(out_7177),
            .b(out_7178),
            .outp(out_7179)
        );        
        

        logic [WIDTH-1:0] out_7180;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7180 (
            .a(out_7171),
            .b(out_7179),
            .outp(out_7180)
        );        
        

        logic [WIDTH-1:0] out_7181;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.9875)
        ) inst_7181 (
            .outp(out_7181)
        );
        

        logic [WIDTH-1:0] out_7182;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7182 (
            .a(out_14),
            .b(out_7181),
            .outp(out_7182)
        );        
        

        logic [WIDTH-1:0] out_7183;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7183 (
            .a(out_6880),
            .b(out_7182),
            .outp(out_7183)
        );        
        

        logic [WIDTH-1:0] out_7184;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.7765)
        ) inst_7184 (
            .outp(out_7184)
        );
        

        logic [WIDTH-1:0] out_7185;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7185 (
            .a(out_7184),
            .b(out_260),
            .outp(out_7185)
        );        
        

        logic [WIDTH-1:0] out_7186;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7186 (
            .a(out_7183),
            .b(out_7185),
            .outp(out_7186)
        );        
        

        logic [WIDTH-1:0] out_7187;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.939)
        ) inst_7187 (
            .outp(out_7187)
        );
        

        logic [WIDTH-1:0] out_7188;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7188 (
            .a(out_260),
            .b(out_7187),
            .outp(out_7188)
        );        
        

        logic [WIDTH-1:0] out_7189;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7189 (
            .a(out_7186),
            .b(out_7188),
            .outp(out_7189)
        );        
        

        logic [WIDTH-1:0] out_7190;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.985)
        ) inst_7190 (
            .outp(out_7190)
        );
        

        logic [WIDTH-1:0] out_7191;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7191 (
            .a(out_7190),
            .b(out_14),
            .outp(out_7191)
        );        
        

        logic [WIDTH-1:0] out_7192;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7192 (
            .in(out_7191),
            .outp(out_7192)
        );
        

        logic [WIDTH-1:0] out_7193;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.84933)
        ) inst_7193 (
            .outp(out_7193)
        );
        

        logic [WIDTH-1:0] out_7194;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7194 (
            .a(out_7193),
            .b(out_241),
            .outp(out_7194)
        );        
        

        logic [WIDTH-1:0] out_7195;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7195 (
            .in(out_7194),
            .outp(out_7195)
        );
        

        logic [WIDTH-1:0] out_7196;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7196 (
            .a(out_7192),
            .b(out_7195),
            .outp(out_7196)
        );        
        

        logic [WIDTH-1:0] out_7197;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7197 (
            .in(out_7196),
            .outp(out_7197)
        );
        

        logic [WIDTH-1:0] out_7198;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7198 (
            .a(out_7197),
            .b(out_250),
            .outp(out_7198)
        );        
        

        logic [WIDTH-1:0] out_7199;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7199 (
            .a(out_7189),
            .b(out_7198),
            .outp(out_7199)
        );        
        

        logic [WIDTH-1:0] out_7200;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7200 (
            .in(out_7199),
            .outp(out_7200)
        );
        

        logic [WIDTH-1:0] out_7201;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7201 (
            .a(out_7181),
            .b(out_14),
            .outp(out_7201)
        );        
        

        logic [WIDTH-1:0] out_7202;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7202 (
            .in(out_7201),
            .outp(out_7202)
        );
        

        logic [WIDTH-1:0] out_7203;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7203 (
            .in(out_7185),
            .outp(out_7203)
        );
        

        logic [WIDTH-1:0] out_7204;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7204 (
            .a(out_7202),
            .b(out_7203),
            .outp(out_7204)
        );        
        

        logic [WIDTH-1:0] out_7205;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7205 (
            .in(out_7204),
            .outp(out_7205)
        );
        

        logic [WIDTH-1:0] out_7206;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7206 (
            .a(out_7205),
            .b(out_275),
            .outp(out_7206)
        );        
        

        logic [WIDTH-1:0] out_7207;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7207 (
            .a(out_7200),
            .b(out_7206),
            .outp(out_7207)
        );        
        

        logic [WIDTH-1:0] out_7208;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7208 (
            .a(out_7180),
            .b(out_7207),
            .outp(out_7208)
        );        
        

        logic [WIDTH-1:0] out_7209;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.925)
        ) inst_7209 (
            .outp(out_7209)
        );
        

        logic [WIDTH-1:0] out_7210;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7210 (
            .a(out_14),
            .b(out_7209),
            .outp(out_7210)
        );        
        

        logic [WIDTH-1:0] out_7211;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.7625)
        ) inst_7211 (
            .outp(out_7211)
        );
        

        logic [WIDTH-1:0] out_7212;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7212 (
            .a(out_7211),
            .b(out_14),
            .outp(out_7212)
        );        
        

        logic [WIDTH-1:0] out_7213;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7213 (
            .a(out_7210),
            .b(out_7212),
            .outp(out_7213)
        );        
        

        logic [WIDTH-1:0] out_7214;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.7765)
        ) inst_7214 (
            .outp(out_7214)
        );
        

        logic [WIDTH-1:0] out_7215;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7215 (
            .a(out_260),
            .b(out_7214),
            .outp(out_7215)
        );        
        

        logic [WIDTH-1:0] out_7216;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7216 (
            .a(out_7213),
            .b(out_7215),
            .outp(out_7216)
        );        
        

        logic [WIDTH-1:0] out_7217;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.614)
        ) inst_7217 (
            .outp(out_7217)
        );
        

        logic [WIDTH-1:0] out_7218;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7218 (
            .a(out_7217),
            .b(out_260),
            .outp(out_7218)
        );        
        

        logic [WIDTH-1:0] out_7219;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7219 (
            .a(out_7216),
            .b(out_7218),
            .outp(out_7219)
        );        
        

        logic [WIDTH-1:0] out_7220;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.765)
        ) inst_7220 (
            .outp(out_7220)
        );
        

        logic [WIDTH-1:0] out_7221;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7221 (
            .a(out_14),
            .b(out_7220),
            .outp(out_7221)
        );        
        

        logic [WIDTH-1:0] out_7222;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7222 (
            .in(out_7221),
            .outp(out_7222)
        );
        

        logic [WIDTH-1:0] out_7223;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.85267)
        ) inst_7223 (
            .outp(out_7223)
        );
        

        logic [WIDTH-1:0] out_7224;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7224 (
            .a(out_241),
            .b(out_7223),
            .outp(out_7224)
        );        
        

        logic [WIDTH-1:0] out_7225;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7225 (
            .in(out_7224),
            .outp(out_7225)
        );
        

        logic [WIDTH-1:0] out_7226;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7226 (
            .a(out_7222),
            .b(out_7225),
            .outp(out_7226)
        );        
        

        logic [WIDTH-1:0] out_7227;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7227 (
            .in(out_7226),
            .outp(out_7227)
        );
        

        logic [WIDTH-1:0] out_7228;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7228 (
            .a(out_7227),
            .b(out_250),
            .outp(out_7228)
        );        
        

        logic [WIDTH-1:0] out_7229;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7229 (
            .a(out_7219),
            .b(out_7228),
            .outp(out_7229)
        );        
        

        logic [WIDTH-1:0] out_7230;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7230 (
            .in(out_7229),
            .outp(out_7230)
        );
        

        logic [WIDTH-1:0] out_7231;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7231 (
            .a(out_14),
            .b(out_7211),
            .outp(out_7231)
        );        
        

        logic [WIDTH-1:0] out_7232;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7232 (
            .in(out_7231),
            .outp(out_7232)
        );
        

        logic [WIDTH-1:0] out_7233;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7233 (
            .in(out_7215),
            .outp(out_7233)
        );
        

        logic [WIDTH-1:0] out_7234;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7234 (
            .a(out_7232),
            .b(out_7233),
            .outp(out_7234)
        );        
        

        logic [WIDTH-1:0] out_7235;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7235 (
            .in(out_7234),
            .outp(out_7235)
        );
        

        logic [WIDTH-1:0] out_7236;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7236 (
            .a(out_7235),
            .b(out_275),
            .outp(out_7236)
        );        
        

        logic [WIDTH-1:0] out_7237;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7237 (
            .a(out_7230),
            .b(out_7236),
            .outp(out_7237)
        );        
        

        logic [WIDTH-1:0] out_7238;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7238 (
            .a(out_7208),
            .b(out_7237),
            .outp(out_7238)
        );        
        

        logic [WIDTH-1:0] out_7239;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.021)
        ) inst_7239 (
            .outp(out_7239)
        );
        

        logic [WIDTH-1:0] out_7240;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7240 (
            .a(out_7239),
            .b(out_3),
            .outp(out_7240)
        );        
        

        logic [WIDTH-1:0] out_7241;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7241 (
            .a(out_7065),
            .b(out_7240),
            .outp(out_7241)
        );        
        

        logic [WIDTH-1:0] out_7242;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.121)
        ) inst_7242 (
            .outp(out_7242)
        );
        

        logic [WIDTH-1:0] out_7243;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7243 (
            .a(out_3),
            .b(out_7242),
            .outp(out_7243)
        );        
        

        logic [WIDTH-1:0] out_7244;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7244 (
            .a(out_7241),
            .b(out_7243),
            .outp(out_7244)
        );        
        

        logic [WIDTH-1:0] out_7245;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7245 (
            .a(out_7238),
            .b(out_7244),
            .outp(out_7245)
        );        
        

        logic [WIDTH-1:0] out_7246;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.05)
        ) inst_7246 (
            .outp(out_7246)
        );
        

        logic [WIDTH-1:0] out_7247;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7247 (
            .a(out_7246),
            .b(out_14),
            .outp(out_7247)
        );        
        

        logic [WIDTH-1:0] out_7248;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7248 (
            .a(out_7121),
            .b(out_7247),
            .outp(out_7248)
        );        
        

        logic [WIDTH-1:0] out_7249;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7249 (
            .a(out_7248),
            .b(out_7073),
            .outp(out_7249)
        );        
        

        logic [WIDTH-1:0] out_7250;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.021)
        ) inst_7250 (
            .outp(out_7250)
        );
        

        logic [WIDTH-1:0] out_7251;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7251 (
            .a(out_3),
            .b(out_7250),
            .outp(out_7251)
        );        
        

        logic [WIDTH-1:0] out_7252;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7252 (
            .a(out_7249),
            .b(out_7251),
            .outp(out_7252)
        );        
        

        logic [WIDTH-1:0] out_7253;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7253 (
            .a(out_7245),
            .b(out_7252),
            .outp(out_7253)
        );        
        

        logic [WIDTH-1:0] out_7254;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7254 (
            .a(out_6924),
            .b(out_7073),
            .outp(out_7254)
        );        
        

        logic [WIDTH-1:0] out_7255;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7255 (
            .a(out_7254),
            .b(out_7251),
            .outp(out_7255)
        );        
        

        logic [WIDTH-1:0] out_7256;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.7)
        ) inst_7256 (
            .outp(out_7256)
        );
        

        logic [WIDTH-1:0] out_7257;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7257 (
            .a(out_14),
            .b(out_7256),
            .outp(out_7257)
        );        
        

        logic [WIDTH-1:0] out_7258;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7258 (
            .a(out_7255),
            .b(out_7257),
            .outp(out_7258)
        );        
        

        logic [WIDTH-1:0] out_7259;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7259 (
            .a(out_7253),
            .b(out_7258),
            .outp(out_7259)
        );        
        

        logic [WIDTH-1:0] out_7260;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7260 (
            .a(out_6924),
            .b(out_7121),
            .outp(out_7260)
        );        
        

        logic [WIDTH-1:0] out_7261;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.12143)
        ) inst_7261 (
            .outp(out_7261)
        );
        

        logic [WIDTH-1:0] out_7262;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7262 (
            .a(out_7261),
            .b(out_194),
            .outp(out_7262)
        );        
        

        logic [WIDTH-1:0] out_7263;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7263 (
            .a(out_7260),
            .b(out_7262),
            .outp(out_7263)
        );        
        

        logic [WIDTH-1:0] out_7264;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.67143)
        ) inst_7264 (
            .outp(out_7264)
        );
        

        logic [WIDTH-1:0] out_7265;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7265 (
            .a(out_7264),
            .b(out_194),
            .outp(out_7265)
        );        
        

        logic [WIDTH-1:0] out_7266;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7266 (
            .in(out_7265),
            .outp(out_7266)
        );
        

        logic [WIDTH-1:0] out_7267;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7267 (
            .a(out_7263),
            .b(out_7266),
            .outp(out_7267)
        );        
        

        logic [WIDTH-1:0] out_7268;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.40179)
        ) inst_7268 (
            .outp(out_7268)
        );
        

        logic [WIDTH-1:0] out_7269;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7269 (
            .a(out_7268),
            .b(out_204),
            .outp(out_7269)
        );        
        

        logic [WIDTH-1:0] out_7270;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7270 (
            .in(out_7269),
            .outp(out_7270)
        );
        

        logic [WIDTH-1:0] out_7271;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7271 (
            .a(out_7131),
            .b(out_7270),
            .outp(out_7271)
        );        
        

        logic [WIDTH-1:0] out_7272;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7272 (
            .in(out_7271),
            .outp(out_7272)
        );
        

        logic [WIDTH-1:0] out_7273;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7273 (
            .a(out_200),
            .b(out_7272),
            .outp(out_7273)
        );        
        

        logic [WIDTH-1:0] out_7274;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7274 (
            .a(out_7267),
            .b(out_7273),
            .outp(out_7274)
        );        
        

        logic [WIDTH-1:0] out_7275;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7275 (
            .in(out_7262),
            .outp(out_7275)
        );
        

        logic [WIDTH-1:0] out_7276;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7276 (
            .a(out_7131),
            .b(out_7275),
            .outp(out_7276)
        );        
        

        logic [WIDTH-1:0] out_7277;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7277 (
            .in(out_7276),
            .outp(out_7277)
        );
        

        logic [WIDTH-1:0] out_7278;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7278 (
            .a(out_7277),
            .b(out_214),
            .outp(out_7278)
        );        
        

        logic [WIDTH-1:0] out_7279;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7279 (
            .a(out_7274),
            .b(out_7278),
            .outp(out_7279)
        );        
        

        logic [WIDTH-1:0] out_7280;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7280 (
            .a(out_7259),
            .b(out_7279),
            .outp(out_7280)
        );        
        

        logic [WIDTH-1:0] out_7281;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.97)
        ) inst_7281 (
            .outp(out_7281)
        );
        

        logic [WIDTH-1:0] out_7282;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7282 (
            .a(out_7281),
            .b(out_3),
            .outp(out_7282)
        );        
        

        logic [WIDTH-1:0] out_7283;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7283 (
            .a(out_7082),
            .b(out_7282),
            .outp(out_7283)
        );        
        

        logic [WIDTH-1:0] out_7284;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.47)
        ) inst_7284 (
            .outp(out_7284)
        );
        

        logic [WIDTH-1:0] out_7285;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7285 (
            .a(out_7284),
            .b(out_3),
            .outp(out_7285)
        );        
        

        logic [WIDTH-1:0] out_7286;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7286 (
            .in(out_7285),
            .outp(out_7286)
        );
        

        logic [WIDTH-1:0] out_7287;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7287 (
            .a(out_7283),
            .b(out_7286),
            .outp(out_7287)
        );        
        

        logic [WIDTH-1:0] out_7288;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.245)
        ) inst_7288 (
            .outp(out_7288)
        );
        

        logic [WIDTH-1:0] out_7289;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7289 (
            .a(out_7288),
            .b(out_3),
            .outp(out_7289)
        );        
        

        logic [WIDTH-1:0] out_7290;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7290 (
            .in(out_7289),
            .outp(out_7290)
        );
        

        logic [WIDTH-1:0] out_7291;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7291 (
            .a(out_6908),
            .b(out_7290),
            .outp(out_7291)
        );        
        

        logic [WIDTH-1:0] out_7292;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7292 (
            .in(out_7291),
            .outp(out_7292)
        );
        

        logic [WIDTH-1:0] out_7293;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7293 (
            .a(out_7292),
            .b(out_21),
            .outp(out_7293)
        );        
        

        logic [WIDTH-1:0] out_7294;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.068)
        ) inst_7294 (
            .outp(out_7294)
        );
        

        logic [WIDTH-1:0] out_7295;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7295 (
            .a(out_7294),
            .b(out_556),
            .outp(out_7295)
        );        
        

        logic [WIDTH-1:0] out_7296;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7296 (
            .a(out_7295),
            .b(out_559),
            .outp(out_7296)
        );        
        

        logic [WIDTH-1:0] out_7297;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7297 (
            .a(out_6891),
            .b(out_7296),
            .outp(out_7297)
        );        
        

        logic [WIDTH-1:0] out_7298;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.272)
        ) inst_7298 (
            .outp(out_7298)
        );
        

        logic [WIDTH-1:0] out_7299;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7299 (
            .a(out_7298),
            .b(out_2653),
            .outp(out_7299)
        );        
        

        logic [WIDTH-1:0] out_7300;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7300 (
            .a(out_7297),
            .b(out_7299),
            .outp(out_7300)
        );        
        

        logic [WIDTH-1:0] out_7301;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7301 (
            .a(out_2653),
            .b(out_7298),
            .outp(out_7301)
        );        
        

        logic [WIDTH-1:0] out_7302;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7302 (
            .a(out_6902),
            .b(out_7301),
            .outp(out_7302)
        );        
        

        logic [WIDTH-1:0] out_7303;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7303 (
            .a(out_559),
            .b(out_7295),
            .outp(out_7303)
        );        
        

        logic [WIDTH-1:0] out_7304;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7304 (
            .a(out_7302),
            .b(out_7303),
            .outp(out_7304)
        );        
        

        logic [WIDTH-1:0] out_7305;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7305 (
            .a(out_7300),
            .b(out_7304),
            .outp(out_7305)
        );        
        

        logic [WIDTH-1:0] out_7306;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7306 (
            .in(out_7305),
            .outp(out_7306)
        );
        

        logic [WIDTH-1:0] out_7307;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7307 (
            .a(out_7293),
            .b(out_7306),
            .outp(out_7307)
        );        
        

        logic [WIDTH-1:0] out_7308;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7308 (
            .a(out_9),
            .b(out_7292),
            .outp(out_7308)
        );        
        

        logic [WIDTH-1:0] out_7309;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7309 (
            .a(out_7307),
            .b(out_7308),
            .outp(out_7309)
        );        
        

        logic [WIDTH-1:0] out_7310;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7310 (
            .a(out_7287),
            .b(out_7309),
            .outp(out_7310)
        );        
        

        logic [WIDTH-1:0] out_7311;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7311 (
            .a(out_7293),
            .b(out_7310),
            .outp(out_7311)
        );        
        

        logic [WIDTH-1:0] out_7312;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7312 (
            .a(out_7280),
            .b(out_7311),
            .outp(out_7312)
        );        
        

        logic [WIDTH-1:0] out_7313;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.36)
        ) inst_7313 (
            .outp(out_7313)
        );
        

        logic [WIDTH-1:0] out_7314;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7314 (
            .a(out_7313),
            .b(out_152),
            .outp(out_7314)
        );        
        

        logic [WIDTH-1:0] out_7315;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.4785)
        ) inst_7315 (
            .outp(out_7315)
        );
        

        logic [WIDTH-1:0] out_7316;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7316 (
            .a(out_7315),
            .b(out_127),
            .outp(out_7316)
        );        
        

        logic [WIDTH-1:0] out_7317;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7317 (
            .a(out_7316),
            .b(out_131),
            .outp(out_7317)
        );        
        

        logic [WIDTH-1:0] out_7318;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7318 (
            .a(out_7314),
            .b(out_7317),
            .outp(out_7318)
        );        
        

        logic [WIDTH-1:0] out_7319;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8935)
        ) inst_7319 (
            .outp(out_7319)
        );
        

        logic [WIDTH-1:0] out_7320;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7320 (
            .a(out_7319),
            .b(out_127),
            .outp(out_7320)
        );        
        

        logic [WIDTH-1:0] out_7321;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7321 (
            .a(out_124),
            .b(out_7320),
            .outp(out_7321)
        );        
        

        logic [WIDTH-1:0] out_7322;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7322 (
            .a(out_7318),
            .b(out_7321),
            .outp(out_7322)
        );        
        

        logic [WIDTH-1:0] out_7323;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7323 (
            .a(out_7312),
            .b(out_7322),
            .outp(out_7323)
        );        
        

        logic [WIDTH-1:0] out_7324;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7324 (
            .a(out_7320),
            .b(out_124),
            .outp(out_7324)
        );        
        

        logic [WIDTH-1:0] out_7325;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7325 (
            .a(out_131),
            .b(out_7316),
            .outp(out_7325)
        );        
        

        logic [WIDTH-1:0] out_7326;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7326 (
            .a(out_7324),
            .b(out_7325),
            .outp(out_7326)
        );        
        

        logic [WIDTH-1:0] out_7327;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7327 (
            .a(out_152),
            .b(out_7313),
            .outp(out_7327)
        );        
        

        logic [WIDTH-1:0] out_7328;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7328 (
            .a(out_7326),
            .b(out_7327),
            .outp(out_7328)
        );        
        

        logic [WIDTH-1:0] out_7329;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7329 (
            .a(out_7323),
            .b(out_7328),
            .outp(out_7329)
        );        
        

        logic [WIDTH-1:0] out_7330;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.415)
        ) inst_7330 (
            .outp(out_7330)
        );
        

        logic [WIDTH-1:0] out_7331;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7331 (
            .a(out_137),
            .b(out_7330),
            .outp(out_7331)
        );        
        

        logic [WIDTH-1:0] out_7332;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7332 (
            .a(out_7324),
            .b(out_7331),
            .outp(out_7332)
        );        
        

        logic [WIDTH-1:0] out_7333;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.5335)
        ) inst_7333 (
            .outp(out_7333)
        );
        

        logic [WIDTH-1:0] out_7334;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7334 (
            .a(out_7333),
            .b(out_127),
            .outp(out_7334)
        );        
        

        logic [WIDTH-1:0] out_7335;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7335 (
            .a(out_131),
            .b(out_7334),
            .outp(out_7335)
        );        
        

        logic [WIDTH-1:0] out_7336;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7336 (
            .a(out_7332),
            .b(out_7335),
            .outp(out_7336)
        );        
        

        logic [WIDTH-1:0] out_7337;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7337 (
            .a(out_7329),
            .b(out_7336),
            .outp(out_7337)
        );        
        

        logic [WIDTH-1:0] out_7338;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7338 (
            .a(out_7334),
            .b(out_131),
            .outp(out_7338)
        );        
        

        logic [WIDTH-1:0] out_7339;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7339 (
            .a(out_7321),
            .b(out_7338),
            .outp(out_7339)
        );        
        

        logic [WIDTH-1:0] out_7340;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7340 (
            .a(out_7330),
            .b(out_137),
            .outp(out_7340)
        );        
        

        logic [WIDTH-1:0] out_7341;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7341 (
            .a(out_7339),
            .b(out_7340),
            .outp(out_7341)
        );        
        

        logic [WIDTH-1:0] out_7342;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7342 (
            .a(out_7337),
            .b(out_7341),
            .outp(out_7342)
        );        
        

        logic [WIDTH-1:0] out_7343;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.7335)
        ) inst_7343 (
            .outp(out_7343)
        );
        

        logic [WIDTH-1:0] out_7344;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7344 (
            .a(out_7343),
            .b(out_131),
            .outp(out_7344)
        );        
        

        logic [WIDTH-1:0] out_7345;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7345 (
            .a(out_7344),
            .b(out_127),
            .outp(out_7345)
        );        
        

        logic [WIDTH-1:0] out_7346;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7346 (
            .in(out_7345),
            .outp(out_7346)
        );
        

        logic [WIDTH-1:0] out_7347;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7347 (
            .a(out_7314),
            .b(out_7346),
            .outp(out_7347)
        );        
        

        logic [WIDTH-1:0] out_7348;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.318501)
        ) inst_7348 (
            .outp(out_7348)
        );
        

        logic [WIDTH-1:0] out_7349;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7349 (
            .a(out_7348),
            .b(out_124),
            .outp(out_7349)
        );        
        

        logic [WIDTH-1:0] out_7350;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7350 (
            .a(out_7349),
            .b(out_127),
            .outp(out_7350)
        );        
        

        logic [WIDTH-1:0] out_7351;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7351 (
            .a(out_7347),
            .b(out_7350),
            .outp(out_7351)
        );        
        

        logic [WIDTH-1:0] out_7352;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7352 (
            .a(out_7342),
            .b(out_7351),
            .outp(out_7352)
        );        
        

        logic [WIDTH-1:0] out_7353;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7353 (
            .a(out_7327),
            .b(out_7345),
            .outp(out_7353)
        );        
        

        logic [WIDTH-1:0] out_7354;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7354 (
            .in(out_7350),
            .outp(out_7354)
        );
        

        logic [WIDTH-1:0] out_7355;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7355 (
            .a(out_7353),
            .b(out_7354),
            .outp(out_7355)
        );        
        

        logic [WIDTH-1:0] out_7356;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7356 (
            .a(out_7352),
            .b(out_7355),
            .outp(out_7356)
        );        
        

        logic [WIDTH-1:0] out_7357;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7357 (
            .a(out_7331),
            .b(out_7354),
            .outp(out_7357)
        );        
        

        logic [WIDTH-1:0] out_7358;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.6785)
        ) inst_7358 (
            .outp(out_7358)
        );
        

        logic [WIDTH-1:0] out_7359;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7359 (
            .a(out_7358),
            .b(out_131),
            .outp(out_7359)
        );        
        

        logic [WIDTH-1:0] out_7360;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7360 (
            .a(out_7359),
            .b(out_127),
            .outp(out_7360)
        );        
        

        logic [WIDTH-1:0] out_7361;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7361 (
            .a(out_7357),
            .b(out_7360),
            .outp(out_7361)
        );        
        

        logic [WIDTH-1:0] out_7362;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7362 (
            .a(out_7356),
            .b(out_7361),
            .outp(out_7362)
        );        
        

        logic [WIDTH-1:0] out_7363;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7363 (
            .a(out_7340),
            .b(out_7350),
            .outp(out_7363)
        );        
        

        logic [WIDTH-1:0] out_7364;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7364 (
            .in(out_7360),
            .outp(out_7364)
        );
        

        logic [WIDTH-1:0] out_7365;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7365 (
            .a(out_7363),
            .b(out_7364),
            .outp(out_7365)
        );        
        

        logic [WIDTH-1:0] out_7366;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7366 (
            .a(out_7362),
            .b(out_7365),
            .outp(out_7366)
        );        
        

        logic [WIDTH-1:0] out_7367;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.34)
        ) inst_7367 (
            .outp(out_7367)
        );
        

        logic [WIDTH-1:0] out_7368;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7368 (
            .a(out_7367),
            .b(out_3),
            .outp(out_7368)
        );        
        

        logic [WIDTH-1:0] out_7369;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7369 (
            .a(out_6925),
            .b(out_7368),
            .outp(out_7369)
        );        
        

        logic [WIDTH-1:0] out_7370;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.44)
        ) inst_7370 (
            .outp(out_7370)
        );
        

        logic [WIDTH-1:0] out_7371;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7371 (
            .a(out_7370),
            .b(out_3),
            .outp(out_7371)
        );        
        

        logic [WIDTH-1:0] out_7372;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7372 (
            .in(out_7371),
            .outp(out_7372)
        );
        

        logic [WIDTH-1:0] out_7373;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7373 (
            .a(out_7369),
            .b(out_7372),
            .outp(out_7373)
        );        
        

        logic [WIDTH-1:0] out_7374;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7374 (
            .a(out_7366),
            .b(out_7373),
            .outp(out_7374)
        );        
        

        logic [WIDTH-1:0] out_7375;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.875)
        ) inst_7375 (
            .outp(out_7375)
        );
        

        logic [WIDTH-1:0] out_7376;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7376 (
            .a(out_7375),
            .b(out_14),
            .outp(out_7376)
        );        
        

        logic [WIDTH-1:0] out_7377;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.688)
        ) inst_7377 (
            .outp(out_7377)
        );
        

        logic [WIDTH-1:0] out_7378;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7378 (
            .a(out_3),
            .b(out_7377),
            .outp(out_7378)
        );        
        

        logic [WIDTH-1:0] out_7379;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7379 (
            .a(out_7376),
            .b(out_7378),
            .outp(out_7379)
        );        
        

        logic [WIDTH-1:0] out_7380;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.587999)
        ) inst_7380 (
            .outp(out_7380)
        );
        

        logic [WIDTH-1:0] out_7381;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7381 (
            .a(out_7380),
            .b(out_3),
            .outp(out_7381)
        );        
        

        logic [WIDTH-1:0] out_7382;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7382 (
            .a(out_7379),
            .b(out_7381),
            .outp(out_7382)
        );        
        

        logic [WIDTH-1:0] out_7383;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7383 (
            .a(out_7382),
            .b(out_7121),
            .outp(out_7383)
        );        
        

        logic [WIDTH-1:0] out_7384;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7384 (
            .a(out_7374),
            .b(out_7383),
            .outp(out_7384)
        );        
        

        logic [WIDTH-1:0] out_7385;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7385 (
            .a(out_6924),
            .b(out_6907),
            .outp(out_7385)
        );        
        

        logic [WIDTH-1:0] out_7386;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7386 (
            .a(out_7385),
            .b(out_7165),
            .outp(out_7386)
        );        
        

        logic [WIDTH-1:0] out_7387;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7387 (
            .a(out_7386),
            .b(out_7381),
            .outp(out_7387)
        );        
        

        logic [WIDTH-1:0] out_7388;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.862999)
        ) inst_7388 (
            .outp(out_7388)
        );
        

        logic [WIDTH-1:0] out_7389;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7389 (
            .a(out_3),
            .b(out_7388),
            .outp(out_7389)
        );        
        

        logic [WIDTH-1:0] out_7390;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7390 (
            .in(out_7389),
            .outp(out_7390)
        );
        

        logic [WIDTH-1:0] out_7391;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7391 (
            .a(out_6908),
            .b(out_7390),
            .outp(out_7391)
        );        
        

        logic [WIDTH-1:0] out_7392;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7392 (
            .in(out_7391),
            .outp(out_7392)
        );
        

        logic [WIDTH-1:0] out_7393;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7393 (
            .a(out_9),
            .b(out_7392),
            .outp(out_7393)
        );        
        

        logic [WIDTH-1:0] out_7394;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7394 (
            .a(out_7387),
            .b(out_7393),
            .outp(out_7394)
        );        
        

        logic [WIDTH-1:0] out_7395;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7395 (
            .a(out_7392),
            .b(out_21),
            .outp(out_7395)
        );        
        

        logic [WIDTH-1:0] out_7396;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7396 (
            .a(out_7394),
            .b(out_7395),
            .outp(out_7396)
        );        
        

        logic [WIDTH-1:0] out_7397;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7397 (
            .a(out_7384),
            .b(out_7396),
            .outp(out_7397)
        );        
        

        logic [WIDTH-1:0] out_7398;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.225)
        ) inst_7398 (
            .outp(out_7398)
        );
        

        logic [WIDTH-1:0] out_7399;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7399 (
            .a(out_7398),
            .b(out_14),
            .outp(out_7399)
        );        
        

        logic [WIDTH-1:0] out_7400;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7400 (
            .a(out_7121),
            .b(out_7399),
            .outp(out_7400)
        );        
        

        logic [WIDTH-1:0] out_7401;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.487999)
        ) inst_7401 (
            .outp(out_7401)
        );
        

        logic [WIDTH-1:0] out_7402;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7402 (
            .a(out_3),
            .b(out_7401),
            .outp(out_7402)
        );        
        

        logic [WIDTH-1:0] out_7403;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7403 (
            .a(out_7400),
            .b(out_7402),
            .outp(out_7403)
        );        
        

        logic [WIDTH-1:0] out_7404;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.387999)
        ) inst_7404 (
            .outp(out_7404)
        );
        

        logic [WIDTH-1:0] out_7405;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7405 (
            .a(out_7404),
            .b(out_3),
            .outp(out_7405)
        );        
        

        logic [WIDTH-1:0] out_7406;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7406 (
            .a(out_7403),
            .b(out_7405),
            .outp(out_7406)
        );        
        

        logic [WIDTH-1:0] out_7407;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7407 (
            .a(out_7397),
            .b(out_7406),
            .outp(out_7407)
        );        
        

        logic [WIDTH-1:0] out_7408;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.212998)
        ) inst_7408 (
            .outp(out_7408)
        );
        

        logic [WIDTH-1:0] out_7409;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7409 (
            .a(out_3),
            .b(out_7408),
            .outp(out_7409)
        );        
        

        logic [WIDTH-1:0] out_7410;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7410 (
            .in(out_7409),
            .outp(out_7410)
        );
        

        logic [WIDTH-1:0] out_7411;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7411 (
            .a(out_6908),
            .b(out_7410),
            .outp(out_7411)
        );        
        

        logic [WIDTH-1:0] out_7412;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7412 (
            .in(out_7411),
            .outp(out_7412)
        );
        

        logic [WIDTH-1:0] out_7413;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7413 (
            .a(out_9),
            .b(out_7412),
            .outp(out_7413)
        );        
        

        logic [WIDTH-1:0] out_7414;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7414 (
            .a(out_7412),
            .b(out_21),
            .outp(out_7414)
        );        
        

        logic [WIDTH-1:0] out_7415;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7415 (
            .a(out_7413),
            .b(out_7414),
            .outp(out_7415)
        );        
        

        logic [WIDTH-1:0] out_7416;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7416 (
            .a(out_7407),
            .b(out_7415),
            .outp(out_7416)
        );        
        

        logic [WIDTH-1:0] out_7417;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.162001)
        ) inst_7417 (
            .outp(out_7417)
        );
        

        logic [WIDTH-1:0] out_7418;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7418 (
            .a(out_7417),
            .b(out_3),
            .outp(out_7418)
        );        
        

        logic [WIDTH-1:0] out_7419;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7419 (
            .a(out_7082),
            .b(out_7418),
            .outp(out_7419)
        );        
        

        logic [WIDTH-1:0] out_7420;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.662001)
        ) inst_7420 (
            .outp(out_7420)
        );
        

        logic [WIDTH-1:0] out_7421;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7421 (
            .a(out_7420),
            .b(out_3),
            .outp(out_7421)
        );        
        

        logic [WIDTH-1:0] out_7422;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7422 (
            .in(out_7421),
            .outp(out_7422)
        );
        

        logic [WIDTH-1:0] out_7423;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7423 (
            .a(out_7419),
            .b(out_7422),
            .outp(out_7423)
        );        
        

        logic [WIDTH-1:0] out_7424;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.437001)
        ) inst_7424 (
            .outp(out_7424)
        );
        

        logic [WIDTH-1:0] out_7425;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7425 (
            .a(out_7424),
            .b(out_3),
            .outp(out_7425)
        );        
        

        logic [WIDTH-1:0] out_7426;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7426 (
            .in(out_7425),
            .outp(out_7426)
        );
        

        logic [WIDTH-1:0] out_7427;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7427 (
            .a(out_6908),
            .b(out_7426),
            .outp(out_7427)
        );        
        

        logic [WIDTH-1:0] out_7428;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7428 (
            .in(out_7427),
            .outp(out_7428)
        );
        

        logic [WIDTH-1:0] out_7429;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7429 (
            .a(out_7428),
            .b(out_21),
            .outp(out_7429)
        );        
        

        logic [WIDTH-1:0] out_7430;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.5708)
        ) inst_7430 (
            .outp(out_7430)
        );
        

        logic [WIDTH-1:0] out_7431;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7431 (
            .a(out_7430),
            .b(out_556),
            .outp(out_7431)
        );        
        

        logic [WIDTH-1:0] out_7432;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7432 (
            .a(out_7431),
            .b(out_559),
            .outp(out_7432)
        );        
        

        logic [WIDTH-1:0] out_7433;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7433 (
            .a(out_6891),
            .b(out_7432),
            .outp(out_7433)
        );        
        

        logic [WIDTH-1:0] out_7434;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.7692)
        ) inst_7434 (
            .outp(out_7434)
        );
        

        logic [WIDTH-1:0] out_7435;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7435 (
            .a(out_7434),
            .b(out_2653),
            .outp(out_7435)
        );        
        

        logic [WIDTH-1:0] out_7436;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7436 (
            .a(out_7433),
            .b(out_7435),
            .outp(out_7436)
        );        
        

        logic [WIDTH-1:0] out_7437;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7437 (
            .a(out_2653),
            .b(out_7434),
            .outp(out_7437)
        );        
        

        logic [WIDTH-1:0] out_7438;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7438 (
            .a(out_6902),
            .b(out_7437),
            .outp(out_7438)
        );        
        

        logic [WIDTH-1:0] out_7439;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7439 (
            .a(out_559),
            .b(out_7431),
            .outp(out_7439)
        );        
        

        logic [WIDTH-1:0] out_7440;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7440 (
            .a(out_7438),
            .b(out_7439),
            .outp(out_7440)
        );        
        

        logic [WIDTH-1:0] out_7441;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7441 (
            .a(out_7436),
            .b(out_7440),
            .outp(out_7441)
        );        
        

        logic [WIDTH-1:0] out_7442;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7442 (
            .in(out_7441),
            .outp(out_7442)
        );
        

        logic [WIDTH-1:0] out_7443;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7443 (
            .a(out_7429),
            .b(out_7442),
            .outp(out_7443)
        );        
        

        logic [WIDTH-1:0] out_7444;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7444 (
            .a(out_9),
            .b(out_7428),
            .outp(out_7444)
        );        
        

        logic [WIDTH-1:0] out_7445;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7445 (
            .a(out_7443),
            .b(out_7444),
            .outp(out_7445)
        );        
        

        logic [WIDTH-1:0] out_7446;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7446 (
            .a(out_7423),
            .b(out_7445),
            .outp(out_7446)
        );        
        

        logic [WIDTH-1:0] out_7447;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7447 (
            .a(out_7429),
            .b(out_7446),
            .outp(out_7447)
        );        
        

        logic [WIDTH-1:0] out_7448;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7448 (
            .a(out_7416),
            .b(out_7447),
            .outp(out_7448)
        );        
        

        logic [WIDTH-1:0] out_7449;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.07)
        ) inst_7449 (
            .outp(out_7449)
        );
        

        logic [WIDTH-1:0] out_7450;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7450 (
            .a(out_7449),
            .b(out_3),
            .outp(out_7450)
        );        
        

        logic [WIDTH-1:0] out_7451;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7451 (
            .a(out_7260),
            .b(out_7450),
            .outp(out_7451)
        );        
        

        logic [WIDTH-1:0] out_7452;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.17)
        ) inst_7452 (
            .outp(out_7452)
        );
        

        logic [WIDTH-1:0] out_7453;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7453 (
            .a(out_7452),
            .b(out_3),
            .outp(out_7453)
        );        
        

        logic [WIDTH-1:0] out_7454;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7454 (
            .in(out_7453),
            .outp(out_7454)
        );
        

        logic [WIDTH-1:0] out_7455;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7455 (
            .a(out_7451),
            .b(out_7454),
            .outp(out_7455)
        );        
        

        logic [WIDTH-1:0] out_7456;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7456 (
            .a(out_7448),
            .b(out_7455),
            .outp(out_7456)
        );        
        

        logic [WIDTH-1:0] out_7457;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.986526)
        ) inst_7457 (
            .outp(out_7457)
        );
        

        logic [WIDTH-1:0] out_7458;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7458 (
            .a(out_7457),
            .b(out_559),
            .outp(out_7458)
        );        
        

        logic [WIDTH-1:0] out_7459;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7459 (
            .a(out_556),
            .b(out_7458),
            .outp(out_7459)
        );        
        

        logic [WIDTH-1:0] out_7460;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7460 (
            .a(out_6360),
            .b(out_7459),
            .outp(out_7460)
        );        
        

        logic [WIDTH-1:0] out_7461;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.04153)
        ) inst_7461 (
            .outp(out_7461)
        );
        

        logic [WIDTH-1:0] out_7462;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7462 (
            .a(out_7461),
            .b(out_2653),
            .outp(out_7462)
        );        
        

        logic [WIDTH-1:0] out_7463;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7463 (
            .a(out_7460),
            .b(out_7462),
            .outp(out_7463)
        );        
        

        logic [WIDTH-1:0] out_7464;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7464 (
            .a(out_2653),
            .b(out_7461),
            .outp(out_7464)
        );        
        

        logic [WIDTH-1:0] out_7465;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7465 (
            .a(out_7458),
            .b(out_556),
            .outp(out_7465)
        );        
        

        logic [WIDTH-1:0] out_7466;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7466 (
            .a(out_7464),
            .b(out_7465),
            .outp(out_7466)
        );        
        

        logic [WIDTH-1:0] out_7467;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7467 (
            .a(out_7466),
            .b(out_6365),
            .outp(out_7467)
        );        
        

        logic [WIDTH-1:0] out_7468;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7468 (
            .a(out_7463),
            .b(out_7467),
            .outp(out_7468)
        );        
        

        logic [WIDTH-1:0] out_7469;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7469 (
            .in(out_7468),
            .outp(out_7469)
        );
        

        logic [WIDTH-1:0] out_7470;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.826)
        ) inst_7470 (
            .outp(out_7470)
        );
        

        logic [WIDTH-1:0] out_7471;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7471 (
            .a(out_3),
            .b(out_7470),
            .outp(out_7471)
        );        
        

        logic [WIDTH-1:0] out_7472;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7472 (
            .in(out_7471),
            .outp(out_7472)
        );
        

        logic [WIDTH-1:0] out_7473;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7473 (
            .a(out_6061),
            .b(out_7472),
            .outp(out_7473)
        );        
        

        logic [WIDTH-1:0] out_7474;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7474 (
            .in(out_7473),
            .outp(out_7474)
        );
        

        logic [WIDTH-1:0] out_7475;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7475 (
            .a(out_9),
            .b(out_7474),
            .outp(out_7475)
        );        
        

        logic [WIDTH-1:0] out_7476;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7476 (
            .a(out_7469),
            .b(out_7475),
            .outp(out_7476)
        );        
        

        logic [WIDTH-1:0] out_7477;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7477 (
            .a(out_7474),
            .b(out_21),
            .outp(out_7477)
        );        
        

        logic [WIDTH-1:0] out_7478;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7478 (
            .a(out_7476),
            .b(out_7477),
            .outp(out_7478)
        );        
        

        logic [WIDTH-1:0] out_7479;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7479 (
            .a(out_6343),
            .b(out_6345),
            .outp(out_7479)
        );        
        

        logic [WIDTH-1:0] out_7480;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.101)
        ) inst_7480 (
            .outp(out_7480)
        );
        

        logic [WIDTH-1:0] out_7481;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7481 (
            .a(out_3),
            .b(out_7480),
            .outp(out_7481)
        );        
        

        logic [WIDTH-1:0] out_7482;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7482 (
            .a(out_7479),
            .b(out_7481),
            .outp(out_7482)
        );        
        

        logic [WIDTH-1:0] out_7483;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.601)
        ) inst_7483 (
            .outp(out_7483)
        );
        

        logic [WIDTH-1:0] out_7484;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7484 (
            .a(out_7483),
            .b(out_3),
            .outp(out_7484)
        );        
        

        logic [WIDTH-1:0] out_7485;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7485 (
            .a(out_7482),
            .b(out_7484),
            .outp(out_7485)
        );        
        

        logic [WIDTH-1:0] out_7486;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7486 (
            .a(out_7478),
            .b(out_7485),
            .outp(out_7486)
        );        
        

        logic [WIDTH-1:0] out_7487;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7487 (
            .a(out_7486),
            .b(out_7477),
            .outp(out_7487)
        );        
        

        logic [WIDTH-1:0] out_7488;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7488 (
            .a(out_7456),
            .b(out_7487),
            .outp(out_7488)
        );        
        

        logic [WIDTH-1:0] out_7489;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.401)
        ) inst_7489 (
            .outp(out_7489)
        );
        

        logic [WIDTH-1:0] out_7490;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7490 (
            .a(out_3),
            .b(out_7489),
            .outp(out_7490)
        );        
        

        logic [WIDTH-1:0] out_7491;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.301)
        ) inst_7491 (
            .outp(out_7491)
        );
        

        logic [WIDTH-1:0] out_7492;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7492 (
            .a(out_7491),
            .b(out_3),
            .outp(out_7492)
        );        
        

        logic [WIDTH-1:0] out_7493;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7493 (
            .a(out_7490),
            .b(out_7492),
            .outp(out_7493)
        );        
        

        logic [WIDTH-1:0] out_7494;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7494 (
            .a(out_7493),
            .b(out_6088),
            .outp(out_7494)
        );        
        

        logic [WIDTH-1:0] out_7495;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7495 (
            .a(out_7494),
            .b(out_6060),
            .outp(out_7495)
        );        
        

        logic [WIDTH-1:0] out_7496;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7496 (
            .a(out_7488),
            .b(out_7495),
            .outp(out_7496)
        );        
        

        logic [WIDTH-1:0] out_7497;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.951)
        ) inst_7497 (
            .outp(out_7497)
        );
        

        logic [WIDTH-1:0] out_7498;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7498 (
            .a(out_3),
            .b(out_7497),
            .outp(out_7498)
        );        
        

        logic [WIDTH-1:0] out_7499;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7499 (
            .a(out_6216),
            .b(out_7498),
            .outp(out_7499)
        );        
        

        logic [WIDTH-1:0] out_7500;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.851)
        ) inst_7500 (
            .outp(out_7500)
        );
        

        logic [WIDTH-1:0] out_7501;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7501 (
            .a(out_7500),
            .b(out_3),
            .outp(out_7501)
        );        
        

        logic [WIDTH-1:0] out_7502;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7502 (
            .a(out_7499),
            .b(out_7501),
            .outp(out_7502)
        );        
        

        logic [WIDTH-1:0] out_7503;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7503 (
            .a(out_7502),
            .b(out_6088),
            .outp(out_7503)
        );        
        

        logic [WIDTH-1:0] out_7504;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7504 (
            .a(out_7496),
            .b(out_7503),
            .outp(out_7504)
        );        
        

        logic [WIDTH-1:0] out_7505;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7505 (
            .a(out_7490),
            .b(out_7501),
            .outp(out_7505)
        );        
        

        logic [WIDTH-1:0] out_7506;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7506 (
            .a(out_7505),
            .b(out_6422),
            .outp(out_7506)
        );        
        

        logic [WIDTH-1:0] out_7507;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.126)
        ) inst_7507 (
            .outp(out_7507)
        );
        

        logic [WIDTH-1:0] out_7508;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7508 (
            .a(out_3),
            .b(out_7507),
            .outp(out_7508)
        );        
        

        logic [WIDTH-1:0] out_7509;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7509 (
            .in(out_7508),
            .outp(out_7509)
        );
        

        logic [WIDTH-1:0] out_7510;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7510 (
            .a(out_7509),
            .b(out_6061),
            .outp(out_7510)
        );        
        

        logic [WIDTH-1:0] out_7511;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7511 (
            .in(out_7510),
            .outp(out_7511)
        );
        

        logic [WIDTH-1:0] out_7512;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7512 (
            .a(out_9),
            .b(out_7511),
            .outp(out_7512)
        );        
        

        logic [WIDTH-1:0] out_7513;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7513 (
            .a(out_7506),
            .b(out_7512),
            .outp(out_7513)
        );        
        

        logic [WIDTH-1:0] out_7514;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7514 (
            .a(out_7511),
            .b(out_21),
            .outp(out_7514)
        );        
        

        logic [WIDTH-1:0] out_7515;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7515 (
            .a(out_7513),
            .b(out_7514),
            .outp(out_7515)
        );        
        

        logic [WIDTH-1:0] out_7516;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7516 (
            .a(out_7515),
            .b(out_6074),
            .outp(out_7516)
        );        
        

        logic [WIDTH-1:0] out_7517;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7517 (
            .a(out_7504),
            .b(out_7516),
            .outp(out_7517)
        );        
        

        logic [WIDTH-1:0] out_7518;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.30055)
        ) inst_7518 (
            .outp(out_7518)
        );
        

        logic [WIDTH-1:0] out_7519;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7519 (
            .a(out_7518),
            .b(out_131),
            .outp(out_7519)
        );        
        

        logic [WIDTH-1:0] out_7520;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7520 (
            .a(out_127),
            .b(out_7519),
            .outp(out_7520)
        );        
        

        logic [WIDTH-1:0] out_7521;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7521 (
            .a(out_6166),
            .b(out_7520),
            .outp(out_7521)
        );        
        

        logic [WIDTH-1:0] out_7522;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(0.775551)
        ) inst_7522 (
            .outp(out_7522)
        );
        

        logic [WIDTH-1:0] out_7523;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7523 (
            .a(out_7522),
            .b(out_124),
            .outp(out_7523)
        );        
        

        logic [WIDTH-1:0] out_7524;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7524 (
            .a(out_7523),
            .b(out_127),
            .outp(out_7524)
        );        
        

        logic [WIDTH-1:0] out_7525;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7525 (
            .a(out_7521),
            .b(out_7524),
            .outp(out_7525)
        );        
        

        logic [WIDTH-1:0] out_7526;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7526 (
            .a(out_7517),
            .b(out_7525),
            .outp(out_7526)
        );        
        

        logic [WIDTH-1:0] out_7527;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7527 (
            .a(out_127),
            .b(out_7523),
            .outp(out_7527)
        );        
        

        logic [WIDTH-1:0] out_7528;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.30055)
        ) inst_7528 (
            .outp(out_7528)
        );
        

        logic [WIDTH-1:0] out_7529;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7529 (
            .a(out_7528),
            .b(out_131),
            .outp(out_7529)
        );        
        

        logic [WIDTH-1:0] out_7530;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7530 (
            .a(out_7529),
            .b(out_127),
            .outp(out_7530)
        );        
        

        logic [WIDTH-1:0] out_7531;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7531 (
            .a(out_7527),
            .b(out_7530),
            .outp(out_7531)
        );        
        

        logic [WIDTH-1:0] out_7532;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7532 (
            .a(out_7531),
            .b(out_6172),
            .outp(out_7532)
        );        
        

        logic [WIDTH-1:0] out_7533;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7533 (
            .a(out_7526),
            .b(out_7532),
            .outp(out_7533)
        );        
        

        logic [WIDTH-1:0] out_7534;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7534 (
            .a(out_7527),
            .b(out_6179),
            .outp(out_7534)
        );        
        

        logic [WIDTH-1:0] out_7535;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.24555)
        ) inst_7535 (
            .outp(out_7535)
        );
        

        logic [WIDTH-1:0] out_7536;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7536 (
            .a(out_7535),
            .b(out_131),
            .outp(out_7536)
        );        
        

        logic [WIDTH-1:0] out_7537;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7537 (
            .a(out_7536),
            .b(out_127),
            .outp(out_7537)
        );        
        

        logic [WIDTH-1:0] out_7538;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7538 (
            .a(out_7534),
            .b(out_7537),
            .outp(out_7538)
        );        
        

        logic [WIDTH-1:0] out_7539;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7539 (
            .a(out_7533),
            .b(out_7538),
            .outp(out_7539)
        );        
        

        logic [WIDTH-1:0] out_7540;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.24555)
        ) inst_7540 (
            .outp(out_7540)
        );
        

        logic [WIDTH-1:0] out_7541;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7541 (
            .a(out_7540),
            .b(out_131),
            .outp(out_7541)
        );        
        

        logic [WIDTH-1:0] out_7542;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7542 (
            .a(out_127),
            .b(out_7541),
            .outp(out_7542)
        );        
        

        logic [WIDTH-1:0] out_7543;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7543 (
            .a(out_7524),
            .b(out_7542),
            .outp(out_7543)
        );        
        

        logic [WIDTH-1:0] out_7544;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7544 (
            .a(out_7543),
            .b(out_6150),
            .outp(out_7544)
        );        
        

        logic [WIDTH-1:0] out_7545;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7545 (
            .a(out_7539),
            .b(out_7544),
            .outp(out_7545)
        );        
        

        logic [WIDTH-1:0] out_7546;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.59555)
        ) inst_7546 (
            .outp(out_7546)
        );
        

        logic [WIDTH-1:0] out_7547;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7547 (
            .a(out_7546),
            .b(out_4477),
            .outp(out_7547)
        );        
        

        logic [WIDTH-1:0] out_7548;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7548 (
            .a(out_6166),
            .b(out_7547),
            .outp(out_7548)
        );        
        

        logic [WIDTH-1:0] out_7549;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7549 (
            .a(out_7548),
            .b(out_6152),
            .outp(out_7549)
        );        
        

        logic [WIDTH-1:0] out_7550;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7550 (
            .a(out_7545),
            .b(out_7549),
            .outp(out_7550)
        );        
        

        logic [WIDTH-1:0] out_7551;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7551 (
            .a(out_6151),
            .b(out_4480),
            .outp(out_7551)
        );        
        

        logic [WIDTH-1:0] out_7552;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7552 (
            .a(out_6172),
            .b(out_7551),
            .outp(out_7552)
        );        
        

        logic [WIDTH-1:0] out_7553;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7553 (
            .a(out_4477),
            .b(out_7546),
            .outp(out_7553)
        );        
        

        logic [WIDTH-1:0] out_7554;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7554 (
            .a(out_7552),
            .b(out_7553),
            .outp(out_7554)
        );        
        

        logic [WIDTH-1:0] out_7555;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7555 (
            .a(out_7550),
            .b(out_7554),
            .outp(out_7555)
        );        
        

        logic [WIDTH-1:0] out_7556;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7556 (
            .a(out_6179),
            .b(out_7551),
            .outp(out_7556)
        );        
        

        logic [WIDTH-1:0] out_7557;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7557 (
            .a(out_4477),
            .b(out_6154),
            .outp(out_7557)
        );        
        

        logic [WIDTH-1:0] out_7558;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7558 (
            .a(out_7556),
            .b(out_7557),
            .outp(out_7558)
        );        
        

        logic [WIDTH-1:0] out_7559;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7559 (
            .a(out_7555),
            .b(out_7558),
            .outp(out_7559)
        );        
        

        logic [WIDTH-1:0] out_7560;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.72857)
        ) inst_7560 (
            .outp(out_7560)
        );
        

        logic [WIDTH-1:0] out_7561;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7561 (
            .a(out_7560),
            .b(out_3),
            .outp(out_7561)
        );        
        

        logic [WIDTH-1:0] out_7562;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7562 (
            .a(out_7561),
            .b(out_1495),
            .outp(out_7562)
        );        
        

        logic [WIDTH-1:0] out_7563;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7563 (
            .in(out_7562),
            .outp(out_7563)
        );
        

        logic [WIDTH-1:0] out_7564;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7564 (
            .a(out_6908),
            .b(out_7563),
            .outp(out_7564)
        );        
        

        logic [WIDTH-1:0] out_7565;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7565 (
            .in(out_7564),
            .outp(out_7565)
        );
        

        logic [WIDTH-1:0] out_7566;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7566 (
            .a(out_9),
            .b(out_7565),
            .outp(out_7566)
        );        
        

        logic [WIDTH-1:0] out_7567;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7567 (
            .a(out_7565),
            .b(out_21),
            .outp(out_7567)
        );        
        

        logic [WIDTH-1:0] out_7568;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7568 (
            .a(out_7566),
            .b(out_7567),
            .outp(out_7568)
        );        
        

        logic [WIDTH-1:0] out_7569;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7569 (
            .a(out_7559),
            .b(out_7568),
            .outp(out_7569)
        );        
        

        logic [WIDTH-1:0] out_7570;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7570 (
            .a(out_7246),
            .b(out_3),
            .outp(out_7570)
        );        
        

        logic [WIDTH-1:0] out_7571;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7571 (
            .a(out_7385),
            .b(out_7570),
            .outp(out_7571)
        );        
        

        logic [WIDTH-1:0] out_7572;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.15)
        ) inst_7572 (
            .outp(out_7572)
        );
        

        logic [WIDTH-1:0] out_7573;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7573 (
            .a(out_7572),
            .b(out_3),
            .outp(out_7573)
        );        
        

        logic [WIDTH-1:0] out_7574;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7574 (
            .in(out_7573),
            .outp(out_7574)
        );
        

        logic [WIDTH-1:0] out_7575;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7575 (
            .a(out_7571),
            .b(out_7574),
            .outp(out_7575)
        );        
        

        logic [WIDTH-1:0] out_7576;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7576 (
            .a(out_7569),
            .b(out_7575),
            .outp(out_7576)
        );        
        

        logic [WIDTH-1:0] out_7577;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7577 (
            .a(out_56),
            .b(out_60),
            .outp(out_7577)
        );        
        

        logic [WIDTH-1:0] out_7578;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7578 (
            .a(out_7577),
            .b(out_6924),
            .outp(out_7578)
        );        
        

        logic [WIDTH-1:0] out_7579;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7579 (
            .a(out_7578),
            .b(out_6448),
            .outp(out_7579)
        );        
        

        logic [WIDTH-1:0] out_7580;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7580 (
            .a(out_7576),
            .b(out_7579),
            .outp(out_7580)
        );        
        

        logic [WIDTH-1:0] out_7581;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7581 (
            .a(out_60),
            .b(out_7376),
            .outp(out_7581)
        );        
        

        logic [WIDTH-1:0] out_7582;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7582 (
            .a(out_7581),
            .b(out_7121),
            .outp(out_7582)
        );        
        

        logic [WIDTH-1:0] out_7583;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7583 (
            .a(out_7582),
            .b(out_7570),
            .outp(out_7583)
        );        
        

        logic [WIDTH-1:0] out_7584;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7584 (
            .a(out_6439),
            .b(out_3),
            .outp(out_7584)
        );        
        

        logic [WIDTH-1:0] out_7585;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7585 (
            .in(out_7584),
            .outp(out_7585)
        );
        

        logic [WIDTH-1:0] out_7586;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7586 (
            .a(out_6908),
            .b(out_7585),
            .outp(out_7586)
        );        
        

        logic [WIDTH-1:0] out_7587;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7587 (
            .in(out_7586),
            .outp(out_7587)
        );
        

        logic [WIDTH-1:0] out_7588;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7588 (
            .a(out_9),
            .b(out_7587),
            .outp(out_7588)
        );        
        

        logic [WIDTH-1:0] out_7589;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7589 (
            .a(out_7583),
            .b(out_7588),
            .outp(out_7589)
        );        
        

        logic [WIDTH-1:0] out_7590;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7590 (
            .a(out_7587),
            .b(out_21),
            .outp(out_7590)
        );        
        

        logic [WIDTH-1:0] out_7591;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7591 (
            .a(out_7589),
            .b(out_7590),
            .outp(out_7591)
        );        
        

        logic [WIDTH-1:0] out_7592;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7592 (
            .a(out_7580),
            .b(out_7591),
            .outp(out_7592)
        );        
        

        logic [WIDTH-1:0] out_7593;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.5)
        ) inst_7593 (
            .outp(out_7593)
        );
        

        logic [WIDTH-1:0] out_7594;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7594 (
            .a(out_7593),
            .b(out_14),
            .outp(out_7594)
        );        
        

        logic [WIDTH-1:0] out_7595;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7595 (
            .a(out_6448),
            .b(out_7594),
            .outp(out_7595)
        );        
        

        logic [WIDTH-1:0] out_7596;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7596 (
            .a(out_6273),
            .b(out_3),
            .outp(out_7596)
        );        
        

        logic [WIDTH-1:0] out_7597;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7597 (
            .a(out_7595),
            .b(out_7596),
            .outp(out_7597)
        );        
        

        logic [WIDTH-1:0] out_7598;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7598 (
            .a(out_6459),
            .b(out_3),
            .outp(out_7598)
        );        
        

        logic [WIDTH-1:0] out_7599;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7599 (
            .in(out_7598),
            .outp(out_7599)
        );
        

        logic [WIDTH-1:0] out_7600;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7600 (
            .a(out_7597),
            .b(out_7599),
            .outp(out_7600)
        );        
        

        logic [WIDTH-1:0] out_7601;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7601 (
            .a(out_7592),
            .b(out_7600),
            .outp(out_7601)
        );        
        

        logic [WIDTH-1:0] out_7602;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7602 (
            .a(out_6924),
            .b(out_7257),
            .outp(out_7602)
        );        
        

        logic [WIDTH-1:0] out_7603;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7603 (
            .a(out_7602),
            .b(out_7596),
            .outp(out_7603)
        );        
        

        logic [WIDTH-1:0] out_7604;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7604 (
            .a(out_7603),
            .b(out_7599),
            .outp(out_7604)
        );        
        

        logic [WIDTH-1:0] out_7605;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7605 (
            .a(out_7601),
            .b(out_7604),
            .outp(out_7605)
        );        
        

        logic [WIDTH-1:0] out_7606;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.6)
        ) inst_7606 (
            .outp(out_7606)
        );
        

        logic [WIDTH-1:0] out_7607;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7607 (
            .a(out_7606),
            .b(out_3),
            .outp(out_7607)
        );        
        

        logic [WIDTH-1:0] out_7608;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7608 (
            .a(out_7065),
            .b(out_7607),
            .outp(out_7608)
        );        
        

        logic [WIDTH-1:0] out_7609;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7609 (
            .a(out_6215),
            .b(out_3),
            .outp(out_7609)
        );        
        

        logic [WIDTH-1:0] out_7610;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7610 (
            .in(out_7609),
            .outp(out_7610)
        );
        

        logic [WIDTH-1:0] out_7611;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7611 (
            .a(out_7608),
            .b(out_7610),
            .outp(out_7611)
        );        
        

        logic [WIDTH-1:0] out_7612;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7612 (
            .a(out_7605),
            .b(out_7611),
            .outp(out_7612)
        );        
        

        logic [WIDTH-1:0] out_7613;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7613 (
            .a(out_6253),
            .b(out_6088),
            .outp(out_7613)
        );        
        

        logic [WIDTH-1:0] out_7614;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.75101)
        ) inst_7614 (
            .outp(out_7614)
        );
        

        logic [WIDTH-1:0] out_7615;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7615 (
            .a(out_3),
            .b(out_7614),
            .outp(out_7615)
        );        
        

        logic [WIDTH-1:0] out_7616;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7616 (
            .a(out_7613),
            .b(out_7615),
            .outp(out_7616)
        );        
        

        logic [WIDTH-1:0] out_7617;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.651)
        ) inst_7617 (
            .outp(out_7617)
        );
        

        logic [WIDTH-1:0] out_7618;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7618 (
            .a(out_7617),
            .b(out_3),
            .outp(out_7618)
        );        
        

        logic [WIDTH-1:0] out_7619;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7619 (
            .a(out_7616),
            .b(out_7618),
            .outp(out_7619)
        );        
        

        logic [WIDTH-1:0] out_7620;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7620 (
            .a(out_7612),
            .b(out_7619),
            .outp(out_7620)
        );        
        

        logic [WIDTH-1:0] out_7621;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7621 (
            .a(out_6088),
            .b(out_6074),
            .outp(out_7621)
        );        
        

        logic [WIDTH-1:0] out_7622;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.30101)
        ) inst_7622 (
            .outp(out_7622)
        );
        

        logic [WIDTH-1:0] out_7623;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7623 (
            .a(out_3),
            .b(out_7622),
            .outp(out_7623)
        );        
        

        logic [WIDTH-1:0] out_7624;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7624 (
            .a(out_7621),
            .b(out_7623),
            .outp(out_7624)
        );        
        

        logic [WIDTH-1:0] out_7625;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.201)
        ) inst_7625 (
            .outp(out_7625)
        );
        

        logic [WIDTH-1:0] out_7626;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7626 (
            .a(out_7625),
            .b(out_3),
            .outp(out_7626)
        );        
        

        logic [WIDTH-1:0] out_7627;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7627 (
            .a(out_7624),
            .b(out_7626),
            .outp(out_7627)
        );        
        

        logic [WIDTH-1:0] out_7628;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7628 (
            .a(out_7620),
            .b(out_7627),
            .outp(out_7628)
        );        
        

        logic [WIDTH-1:0] out_7629;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7629 (
            .a(out_7615),
            .b(out_6074),
            .outp(out_7629)
        );        
        

        logic [WIDTH-1:0] out_7630;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7630 (
            .a(out_7629),
            .b(out_7626),
            .outp(out_7630)
        );        
        

        logic [WIDTH-1:0] out_7631;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7631 (
            .a(out_7630),
            .b(out_6077),
            .outp(out_7631)
        );        
        

        logic [WIDTH-1:0] out_7632;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.476)
        ) inst_7632 (
            .outp(out_7632)
        );
        

        logic [WIDTH-1:0] out_7633;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7633 (
            .a(out_3),
            .b(out_7632),
            .outp(out_7633)
        );        
        

        logic [WIDTH-1:0] out_7634;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7634 (
            .in(out_7633),
            .outp(out_7634)
        );
        

        logic [WIDTH-1:0] out_7635;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7635 (
            .a(out_6061),
            .b(out_7634),
            .outp(out_7635)
        );        
        

        logic [WIDTH-1:0] out_7636;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7636 (
            .in(out_7635),
            .outp(out_7636)
        );
        

        logic [WIDTH-1:0] out_7637;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7637 (
            .a(out_9),
            .b(out_7636),
            .outp(out_7637)
        );        
        

        logic [WIDTH-1:0] out_7638;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7638 (
            .a(out_7631),
            .b(out_7637),
            .outp(out_7638)
        );        
        

        logic [WIDTH-1:0] out_7639;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7639 (
            .a(out_7636),
            .b(out_21),
            .outp(out_7639)
        );        
        

        logic [WIDTH-1:0] out_7640;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7640 (
            .a(out_7638),
            .b(out_7639),
            .outp(out_7640)
        );        
        

        logic [WIDTH-1:0] out_7641;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7641 (
            .a(out_7628),
            .b(out_7640),
            .outp(out_7641)
        );        
        

        logic [WIDTH-1:0] out_7642;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7642 (
            .a(out_6509),
            .b(out_6726),
            .outp(out_7642)
        );        
        

        logic [WIDTH-1:0] out_7643;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7643 (
            .a(out_5145),
            .b(out_3),
            .outp(out_7643)
        );        
        

        logic [WIDTH-1:0] out_7644;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7644 (
            .a(out_7642),
            .b(out_7643),
            .outp(out_7644)
        );        
        

        logic [WIDTH-1:0] out_7645;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7645 (
            .in(out_798),
            .outp(out_7645)
        );
        

        logic [WIDTH-1:0] out_7646;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7646 (
            .a(out_7644),
            .b(out_7645),
            .outp(out_7646)
        );        
        

        logic [WIDTH-1:0] out_7647;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7647 (
            .in(out_791),
            .outp(out_7647)
        );
        

        logic [WIDTH-1:0] out_7648;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7648 (
            .a(out_6498),
            .b(out_7647),
            .outp(out_7648)
        );        
        

        logic [WIDTH-1:0] out_7649;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7649 (
            .in(out_7648),
            .outp(out_7649)
        );
        

        logic [WIDTH-1:0] out_7650;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7650 (
            .a(out_9),
            .b(out_7649),
            .outp(out_7650)
        );        
        

        logic [WIDTH-1:0] out_7651;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7651 (
            .a(out_7646),
            .b(out_7650),
            .outp(out_7651)
        );        
        

        logic [WIDTH-1:0] out_7652;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7652 (
            .a(out_7649),
            .b(out_21),
            .outp(out_7652)
        );        
        

        logic [WIDTH-1:0] out_7653;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7653 (
            .a(out_7651),
            .b(out_7652),
            .outp(out_7653)
        );        
        

        logic [WIDTH-1:0] out_7654;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7654 (
            .a(out_7641),
            .b(out_7653),
            .outp(out_7654)
        );        
        

        logic [WIDTH-1:0] out_7655;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7655 (
            .a(out_6655),
            .b(out_14),
            .outp(out_7655)
        );        
        

        logic [WIDTH-1:0] out_7656;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7656 (
            .a(out_6477),
            .b(out_7655),
            .outp(out_7656)
        );        
        

        logic [WIDTH-1:0] out_7657;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7657 (
            .a(out_2111),
            .b(out_3),
            .outp(out_7657)
        );        
        

        logic [WIDTH-1:0] out_7658;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7658 (
            .a(out_7656),
            .b(out_7657),
            .outp(out_7658)
        );        
        

        logic [WIDTH-1:0] out_7659;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7659 (
            .a(out_7209),
            .b(out_3),
            .outp(out_7659)
        );        
        

        logic [WIDTH-1:0] out_7660;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7660 (
            .in(out_7659),
            .outp(out_7660)
        );
        

        logic [WIDTH-1:0] out_7661;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7661 (
            .a(out_7658),
            .b(out_7660),
            .outp(out_7661)
        );        
        

        logic [WIDTH-1:0] out_7662;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7662 (
            .a(out_7654),
            .b(out_7661),
            .outp(out_7662)
        );        
        

        logic [WIDTH-1:0] out_7663;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7663 (
            .a(out_3253),
            .b(out_14),
            .outp(out_7663)
        );        
        

        logic [WIDTH-1:0] out_7664;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7664 (
            .a(out_6824),
            .b(out_7663),
            .outp(out_7664)
        );        
        

        logic [WIDTH-1:0] out_7665;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.675)
        ) inst_7665 (
            .outp(out_7665)
        );
        

        logic [WIDTH-1:0] out_7666;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7666 (
            .a(out_7665),
            .b(out_3),
            .outp(out_7666)
        );        
        

        logic [WIDTH-1:0] out_7667;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7667 (
            .a(out_7664),
            .b(out_7666),
            .outp(out_7667)
        );        
        

        logic [WIDTH-1:0] out_7668;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.075)
        ) inst_7668 (
            .outp(out_7668)
        );
        

        logic [WIDTH-1:0] out_7669;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7669 (
            .a(out_7668),
            .b(out_3),
            .outp(out_7669)
        );        
        

        logic [WIDTH-1:0] out_7670;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7670 (
            .in(out_7669),
            .outp(out_7670)
        );
        

        logic [WIDTH-1:0] out_7671;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7671 (
            .a(out_7667),
            .b(out_7670),
            .outp(out_7671)
        );        
        

        logic [WIDTH-1:0] out_7672;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7672 (
            .a(out_7662),
            .b(out_7671),
            .outp(out_7672)
        );        
        

        logic [WIDTH-1:0] out_7673;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7673 (
            .a(out_6462),
            .b(out_7666),
            .outp(out_7673)
        );        
        

        logic [WIDTH-1:0] out_7674;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7674 (
            .a(out_7673),
            .b(out_7670),
            .outp(out_7674)
        );        
        

        logic [WIDTH-1:0] out_7675;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7675 (
            .a(out_14),
            .b(out_6655),
            .outp(out_7675)
        );        
        

        logic [WIDTH-1:0] out_7676;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7676 (
            .a(out_7674),
            .b(out_7675),
            .outp(out_7676)
        );        
        

        logic [WIDTH-1:0] out_7677;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7677 (
            .in(out_7675),
            .outp(out_7677)
        );
        

        logic [WIDTH-1:0] out_7678;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7678 (
            .in(out_7666),
            .outp(out_7678)
        );
        

        logic [WIDTH-1:0] out_7679;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7679 (
            .a(out_7677),
            .b(out_7678),
            .outp(out_7679)
        );        
        

        logic [WIDTH-1:0] out_7680;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7680 (
            .in(out_7679),
            .outp(out_7680)
        );
        

        logic [WIDTH-1:0] out_7681;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7681 (
            .a(out_336),
            .b(out_7680),
            .outp(out_7681)
        );        
        

        logic [WIDTH-1:0] out_7682;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7682 (
            .a(out_7676),
            .b(out_7681),
            .outp(out_7682)
        );        
        

        logic [WIDTH-1:0] out_7683;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7683 (
            .a(out_7680),
            .b(out_343),
            .outp(out_7683)
        );        
        

        logic [WIDTH-1:0] out_7684;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7684 (
            .a(out_7682),
            .b(out_7683),
            .outp(out_7684)
        );        
        

        logic [WIDTH-1:0] out_7685;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7685 (
            .a(out_7672),
            .b(out_7684),
            .outp(out_7685)
        );        
        

        logic [WIDTH-1:0] out_7686;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7686 (
            .a(out_6076),
            .b(out_3),
            .outp(out_7686)
        );        
        

        logic [WIDTH-1:0] out_7687;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7687 (
            .a(out_7656),
            .b(out_7686),
            .outp(out_7687)
        );        
        

        logic [WIDTH-1:0] out_7688;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.125)
        ) inst_7688 (
            .outp(out_7688)
        );
        

        logic [WIDTH-1:0] out_7689;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7689 (
            .a(out_7688),
            .b(out_3),
            .outp(out_7689)
        );        
        

        logic [WIDTH-1:0] out_7690;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7690 (
            .in(out_7689),
            .outp(out_7690)
        );
        

        logic [WIDTH-1:0] out_7691;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7691 (
            .a(out_7687),
            .b(out_7690),
            .outp(out_7691)
        );        
        

        logic [WIDTH-1:0] out_7692;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7692 (
            .a(out_7685),
            .b(out_7691),
            .outp(out_7692)
        );        
        

        logic [WIDTH-1:0] out_7693;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(4.875)
        ) inst_7693 (
            .outp(out_7693)
        );
        

        logic [WIDTH-1:0] out_7694;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7694 (
            .a(out_7693),
            .b(out_3),
            .outp(out_7694)
        );        
        

        logic [WIDTH-1:0] out_7695;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7695 (
            .a(out_7664),
            .b(out_7694),
            .outp(out_7695)
        );        
        

        logic [WIDTH-1:0] out_7696;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7696 (
            .in(out_5283),
            .outp(out_7696)
        );
        

        logic [WIDTH-1:0] out_7697;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7697 (
            .a(out_7695),
            .b(out_7696),
            .outp(out_7697)
        );        
        

        logic [WIDTH-1:0] out_7698;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7698 (
            .a(out_7692),
            .b(out_7697),
            .outp(out_7698)
        );        
        

        logic [WIDTH-1:0] out_7699;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7699 (
            .a(out_6462),
            .b(out_7675),
            .outp(out_7699)
        );        
        

        logic [WIDTH-1:0] out_7700;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7700 (
            .a(out_7699),
            .b(out_7694),
            .outp(out_7700)
        );        
        

        logic [WIDTH-1:0] out_7701;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7701 (
            .a(out_7700),
            .b(out_7696),
            .outp(out_7701)
        );        
        

        logic [WIDTH-1:0] out_7702;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7702 (
            .in(out_7694),
            .outp(out_7702)
        );
        

        logic [WIDTH-1:0] out_7703;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7703 (
            .a(out_7677),
            .b(out_7702),
            .outp(out_7703)
        );        
        

        logic [WIDTH-1:0] out_7704;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7704 (
            .in(out_7703),
            .outp(out_7704)
        );
        

        logic [WIDTH-1:0] out_7705;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7705 (
            .a(out_336),
            .b(out_7704),
            .outp(out_7705)
        );        
        

        logic [WIDTH-1:0] out_7706;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7706 (
            .a(out_7701),
            .b(out_7705),
            .outp(out_7706)
        );        
        

        logic [WIDTH-1:0] out_7707;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7707 (
            .a(out_7704),
            .b(out_343),
            .outp(out_7707)
        );        
        

        logic [WIDTH-1:0] out_7708;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7708 (
            .a(out_7706),
            .b(out_7707),
            .outp(out_7708)
        );        
        

        logic [WIDTH-1:0] out_7709;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7709 (
            .a(out_7698),
            .b(out_7708),
            .outp(out_7709)
        );        
        

        logic [WIDTH-1:0] out_7710;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7710 (
            .a(out_5286),
            .b(out_6462),
            .outp(out_7710)
        );        
        

        logic [WIDTH-1:0] out_7711;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7711 (
            .a(out_7710),
            .b(out_6509),
            .outp(out_7711)
        );        
        

        logic [WIDTH-1:0] out_7712;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.475)
        ) inst_7712 (
            .outp(out_7712)
        );
        

        logic [WIDTH-1:0] out_7713;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7713 (
            .a(out_7712),
            .b(out_3),
            .outp(out_7713)
        );        
        

        logic [WIDTH-1:0] out_7714;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7714 (
            .in(out_7713),
            .outp(out_7714)
        );
        

        logic [WIDTH-1:0] out_7715;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7715 (
            .a(out_7711),
            .b(out_7714),
            .outp(out_7715)
        );        
        

        logic [WIDTH-1:0] out_7716;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7716 (
            .a(out_7709),
            .b(out_7715),
            .outp(out_7716)
        );        
        

        logic [WIDTH-1:0] out_7717;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.825)
        ) inst_7717 (
            .outp(out_7717)
        );
        

        logic [WIDTH-1:0] out_7718;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7718 (
            .a(out_7717),
            .b(out_3),
            .outp(out_7718)
        );        
        

        logic [WIDTH-1:0] out_7719;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7719 (
            .a(out_7642),
            .b(out_7718),
            .outp(out_7719)
        );        
        

        logic [WIDTH-1:0] out_7720;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.925)
        ) inst_7720 (
            .outp(out_7720)
        );
        

        logic [WIDTH-1:0] out_7721;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7721 (
            .a(out_7720),
            .b(out_3),
            .outp(out_7721)
        );        
        

        logic [WIDTH-1:0] out_7722;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7722 (
            .in(out_7721),
            .outp(out_7722)
        );
        

        logic [WIDTH-1:0] out_7723;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7723 (
            .a(out_7719),
            .b(out_7722),
            .outp(out_7723)
        );        
        

        logic [WIDTH-1:0] out_7724;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7724 (
            .a(out_7716),
            .b(out_7723),
            .outp(out_7724)
        );        
        

        logic [WIDTH-1:0] out_7725;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7725 (
            .a(out_7710),
            .b(out_6497),
            .outp(out_7725)
        );        
        

        logic [WIDTH-1:0] out_7726;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7726 (
            .a(out_7725),
            .b(out_7722),
            .outp(out_7726)
        );        
        

        logic [WIDTH-1:0] out_7727;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.65)
        ) inst_7727 (
            .outp(out_7727)
        );
        

        logic [WIDTH-1:0] out_7728;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7728 (
            .a(out_7727),
            .b(out_3),
            .outp(out_7728)
        );        
        

        logic [WIDTH-1:0] out_7729;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7729 (
            .in(out_7728),
            .outp(out_7729)
        );
        

        logic [WIDTH-1:0] out_7730;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7730 (
            .a(out_6498),
            .b(out_7729),
            .outp(out_7730)
        );        
        

        logic [WIDTH-1:0] out_7731;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7731 (
            .in(out_7730),
            .outp(out_7731)
        );
        

        logic [WIDTH-1:0] out_7732;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7732 (
            .a(out_9),
            .b(out_7731),
            .outp(out_7732)
        );        
        

        logic [WIDTH-1:0] out_7733;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7733 (
            .a(out_7726),
            .b(out_7732),
            .outp(out_7733)
        );        
        

        logic [WIDTH-1:0] out_7734;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7734 (
            .a(out_7731),
            .b(out_21),
            .outp(out_7734)
        );        
        

        logic [WIDTH-1:0] out_7735;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7735 (
            .a(out_7733),
            .b(out_7734),
            .outp(out_7735)
        );        
        

        logic [WIDTH-1:0] out_7736;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7736 (
            .a(out_7724),
            .b(out_7735),
            .outp(out_7736)
        );        
        

        logic [WIDTH-1:0] out_7737;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7737 (
            .a(out_6664),
            .b(out_6462),
            .outp(out_7737)
        );        
        

        logic [WIDTH-1:0] out_7738;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7738 (
            .a(out_7737),
            .b(out_6477),
            .outp(out_7738)
        );        
        

        logic [WIDTH-1:0] out_7739;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7739 (
            .a(out_7736),
            .b(out_7738),
            .outp(out_7739)
        );        
        

        logic [WIDTH-1:0] out_7740;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7740 (
            .a(out_4167),
            .b(out_6477),
            .outp(out_7740)
        );        
        

        logic [WIDTH-1:0] out_7741;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7741 (
            .a(out_7740),
            .b(out_6679),
            .outp(out_7741)
        );        
        

        logic [WIDTH-1:0] out_7742;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.3)
        ) inst_7742 (
            .outp(out_7742)
        );
        

        logic [WIDTH-1:0] out_7743;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7743 (
            .a(out_7742),
            .b(out_3),
            .outp(out_7743)
        );        
        

        logic [WIDTH-1:0] out_7744;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7744 (
            .a(out_7741),
            .b(out_7743),
            .outp(out_7744)
        );        
        

        logic [WIDTH-1:0] out_7745;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7745 (
            .a(out_7739),
            .b(out_7744),
            .outp(out_7745)
        );        
        

        logic [WIDTH-1:0] out_7746;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7746 (
            .a(out_4167),
            .b(out_6509),
            .outp(out_7746)
        );        
        

        logic [WIDTH-1:0] out_7747;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7747 (
            .a(out_7746),
            .b(out_7743),
            .outp(out_7747)
        );        
        

        logic [WIDTH-1:0] out_7748;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7748 (
            .a(out_3040),
            .b(out_14),
            .outp(out_7748)
        );        
        

        logic [WIDTH-1:0] out_7749;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7749 (
            .a(out_7747),
            .b(out_7748),
            .outp(out_7749)
        );        
        

        logic [WIDTH-1:0] out_7750;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7750 (
            .a(out_7745),
            .b(out_7749),
            .outp(out_7750)
        );        
        

        logic [WIDTH-1:0] out_7751;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7751 (
            .a(out_4167),
            .b(out_6460),
            .outp(out_7751)
        );        
        

        logic [WIDTH-1:0] out_7752;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7752 (
            .a(out_7751),
            .b(out_6462),
            .outp(out_7752)
        );        
        

        logic [WIDTH-1:0] out_7753;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7753 (
            .a(out_7752),
            .b(out_7743),
            .outp(out_7753)
        );        
        

        logic [WIDTH-1:0] out_7754;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7754 (
            .a(out_7750),
            .b(out_7753),
            .outp(out_7754)
        );        
        

        logic [WIDTH-1:0] out_7755;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.025)
        ) inst_7755 (
            .outp(out_7755)
        );
        

        logic [WIDTH-1:0] out_7756;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7756 (
            .a(out_7755),
            .b(out_14),
            .outp(out_7756)
        );        
        

        logic [WIDTH-1:0] out_7757;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.1875)
        ) inst_7757 (
            .outp(out_7757)
        );
        

        logic [WIDTH-1:0] out_7758;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7758 (
            .a(out_14),
            .b(out_7757),
            .outp(out_7758)
        );        
        

        logic [WIDTH-1:0] out_7759;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7759 (
            .a(out_7756),
            .b(out_7758),
            .outp(out_7759)
        );        
        

        logic [WIDTH-1:0] out_7760;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5875)
        ) inst_7760 (
            .outp(out_7760)
        );
        

        logic [WIDTH-1:0] out_7761;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7761 (
            .a(out_7760),
            .b(out_260),
            .outp(out_7761)
        );        
        

        logic [WIDTH-1:0] out_7762;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7762 (
            .in(out_7761),
            .outp(out_7762)
        );
        

        logic [WIDTH-1:0] out_7763;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7763 (
            .a(out_7759),
            .b(out_7762),
            .outp(out_7763)
        );        
        

        logic [WIDTH-1:0] out_7764;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.425)
        ) inst_7764 (
            .outp(out_7764)
        );
        

        logic [WIDTH-1:0] out_7765;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7765 (
            .a(out_7764),
            .b(out_260),
            .outp(out_7765)
        );        
        

        logic [WIDTH-1:0] out_7766;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7766 (
            .a(out_7763),
            .b(out_7765),
            .outp(out_7766)
        );        
        

        logic [WIDTH-1:0] out_7767;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.185)
        ) inst_7767 (
            .outp(out_7767)
        );
        

        logic [WIDTH-1:0] out_7768;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7768 (
            .a(out_7767),
            .b(out_14),
            .outp(out_7768)
        );        
        

        logic [WIDTH-1:0] out_7769;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7769 (
            .in(out_7768),
            .outp(out_7769)
        );
        

        logic [WIDTH-1:0] out_7770;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.06)
        ) inst_7770 (
            .outp(out_7770)
        );
        

        logic [WIDTH-1:0] out_7771;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7771 (
            .a(out_7770),
            .b(out_241),
            .outp(out_7771)
        );        
        

        logic [WIDTH-1:0] out_7772;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7772 (
            .in(out_7771),
            .outp(out_7772)
        );
        

        logic [WIDTH-1:0] out_7773;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7773 (
            .in(out_7772),
            .outp(out_7773)
        );
        

        logic [WIDTH-1:0] out_7774;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7774 (
            .a(out_7769),
            .b(out_7773),
            .outp(out_7774)
        );        
        

        logic [WIDTH-1:0] out_7775;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7775 (
            .in(out_7774),
            .outp(out_7775)
        );
        

        logic [WIDTH-1:0] out_7776;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7776 (
            .a(out_7775),
            .b(out_250),
            .outp(out_7776)
        );        
        

        logic [WIDTH-1:0] out_7777;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7777 (
            .a(out_7766),
            .b(out_7776),
            .outp(out_7777)
        );        
        

        logic [WIDTH-1:0] out_7778;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7778 (
            .in(out_7777),
            .outp(out_7778)
        );
        

        logic [WIDTH-1:0] out_7779;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7779 (
            .a(out_7757),
            .b(out_14),
            .outp(out_7779)
        );        
        

        logic [WIDTH-1:0] out_7780;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7780 (
            .in(out_7779),
            .outp(out_7780)
        );
        

        logic [WIDTH-1:0] out_7781;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7781 (
            .in(out_7762),
            .outp(out_7781)
        );
        

        logic [WIDTH-1:0] out_7782;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7782 (
            .a(out_7780),
            .b(out_7781),
            .outp(out_7782)
        );        
        

        logic [WIDTH-1:0] out_7783;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7783 (
            .in(out_7782),
            .outp(out_7783)
        );
        

        logic [WIDTH-1:0] out_7784;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7784 (
            .a(out_7783),
            .b(out_275),
            .outp(out_7784)
        );        
        

        logic [WIDTH-1:0] out_7785;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7785 (
            .a(out_7778),
            .b(out_7784),
            .outp(out_7785)
        );        
        

        logic [WIDTH-1:0] out_7786;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7786 (
            .a(out_7754),
            .b(out_7785),
            .outp(out_7786)
        );        
        

        logic [WIDTH-1:0] out_7787;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.125)
        ) inst_7787 (
            .outp(out_7787)
        );
        

        logic [WIDTH-1:0] out_7788;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7788 (
            .a(out_14),
            .b(out_7787),
            .outp(out_7788)
        );        
        

        logic [WIDTH-1:0] out_7789;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.9625)
        ) inst_7789 (
            .outp(out_7789)
        );
        

        logic [WIDTH-1:0] out_7790;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7790 (
            .a(out_7789),
            .b(out_14),
            .outp(out_7790)
        );        
        

        logic [WIDTH-1:0] out_7791;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7791 (
            .a(out_7788),
            .b(out_7790),
            .outp(out_7791)
        );        
        

        logic [WIDTH-1:0] out_7792;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.5875)
        ) inst_7792 (
            .outp(out_7792)
        );
        

        logic [WIDTH-1:0] out_7793;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7793 (
            .a(out_7792),
            .b(out_260),
            .outp(out_7793)
        );        
        

        logic [WIDTH-1:0] out_7794;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7794 (
            .a(out_7791),
            .b(out_7793),
            .outp(out_7794)
        );        
        

        logic [WIDTH-1:0] out_7795;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.75)
        ) inst_7795 (
            .outp(out_7795)
        );
        

        logic [WIDTH-1:0] out_7796;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7796 (
            .a(out_7795),
            .b(out_260),
            .outp(out_7796)
        );        
        

        logic [WIDTH-1:0] out_7797;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7797 (
            .in(out_7796),
            .outp(out_7797)
        );
        

        logic [WIDTH-1:0] out_7798;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7798 (
            .a(out_7794),
            .b(out_7797),
            .outp(out_7798)
        );        
        

        logic [WIDTH-1:0] out_7799;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(5.965)
        ) inst_7799 (
            .outp(out_7799)
        );
        

        logic [WIDTH-1:0] out_7800;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7800 (
            .a(out_14),
            .b(out_7799),
            .outp(out_7800)
        );        
        

        logic [WIDTH-1:0] out_7801;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7801 (
            .in(out_7800),
            .outp(out_7801)
        );
        

        logic [WIDTH-1:0] out_7802;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(1.05667)
        ) inst_7802 (
            .outp(out_7802)
        );
        

        logic [WIDTH-1:0] out_7803;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7803 (
            .a(out_7802),
            .b(out_241),
            .outp(out_7803)
        );        
        

        logic [WIDTH-1:0] out_7804;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7804 (
            .in(out_7803),
            .outp(out_7804)
        );
        

        logic [WIDTH-1:0] out_7805;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7805 (
            .a(out_7801),
            .b(out_7804),
            .outp(out_7805)
        );        
        

        logic [WIDTH-1:0] out_7806;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7806 (
            .in(out_7805),
            .outp(out_7806)
        );
        

        logic [WIDTH-1:0] out_7807;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7807 (
            .a(out_7806),
            .b(out_250),
            .outp(out_7807)
        );        
        

        logic [WIDTH-1:0] out_7808;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7808 (
            .a(out_7798),
            .b(out_7807),
            .outp(out_7808)
        );        
        

        logic [WIDTH-1:0] out_7809;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7809 (
            .in(out_7808),
            .outp(out_7809)
        );
        

        logic [WIDTH-1:0] out_7810;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7810 (
            .a(out_14),
            .b(out_7789),
            .outp(out_7810)
        );        
        

        logic [WIDTH-1:0] out_7811;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7811 (
            .in(out_7810),
            .outp(out_7811)
        );
        

        logic [WIDTH-1:0] out_7812;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7812 (
            .in(out_7793),
            .outp(out_7812)
        );
        

        logic [WIDTH-1:0] out_7813;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7813 (
            .a(out_7811),
            .b(out_7812),
            .outp(out_7813)
        );        
        

        logic [WIDTH-1:0] out_7814;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7814 (
            .in(out_7813),
            .outp(out_7814)
        );
        

        logic [WIDTH-1:0] out_7815;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7815 (
            .a(out_7814),
            .b(out_275),
            .outp(out_7815)
        );        
        

        logic [WIDTH-1:0] out_7816;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7816 (
            .a(out_7809),
            .b(out_7815),
            .outp(out_7816)
        );        
        

        logic [WIDTH-1:0] out_7817;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7817 (
            .a(out_7786),
            .b(out_7816),
            .outp(out_7817)
        );        
        

        logic [WIDTH-1:0] out_7818;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.75)
        ) inst_7818 (
            .outp(out_7818)
        );
        

        logic [WIDTH-1:0] out_7819;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7819 (
            .a(out_7818),
            .b(out_3),
            .outp(out_7819)
        );        
        

        logic [WIDTH-1:0] out_7820;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7820 (
            .a(out_6510),
            .b(out_7819),
            .outp(out_7820)
        );        
        

        logic [WIDTH-1:0] out_7821;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.85)
        ) inst_7821 (
            .outp(out_7821)
        );
        

        logic [WIDTH-1:0] out_7822;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7822 (
            .a(out_7821),
            .b(out_3),
            .outp(out_7822)
        );        
        

        logic [WIDTH-1:0] out_7823;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7823 (
            .in(out_7822),
            .outp(out_7823)
        );
        

        logic [WIDTH-1:0] out_7824;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7824 (
            .a(out_7820),
            .b(out_7823),
            .outp(out_7824)
        );        
        

        logic [WIDTH-1:0] out_7825;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7825 (
            .a(out_7817),
            .b(out_7824),
            .outp(out_7825)
        );        
        

        logic [WIDTH-1:0] out_7826;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(2.8)
        ) inst_7826 (
            .outp(out_7826)
        );
        

        logic [WIDTH-1:0] out_7827;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7827 (
            .a(out_7826),
            .b(out_3),
            .outp(out_7827)
        );        
        

        logic [WIDTH-1:0] out_7828;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7828 (
            .in(out_7827),
            .outp(out_7828)
        );
        

        logic [WIDTH-1:0] out_7829;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7829 (
            .a(out_6519),
            .b(out_7828),
            .outp(out_7829)
        );        
        

        logic [WIDTH-1:0] out_7830;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7830 (
            .in(out_7829),
            .outp(out_7830)
        );
        

        logic [WIDTH-1:0] out_7831;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7831 (
            .a(out_7830),
            .b(out_460),
            .outp(out_7831)
        );        
        

        logic [WIDTH-1:0] out_7832;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7832 (
            .a(out_7825),
            .b(out_7831),
            .outp(out_7832)
        );        
        

        logic [WIDTH-1:0] out_7833;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7833 (
            .a(out_6729),
            .b(out_7643),
            .outp(out_7833)
        );        
        

        logic [WIDTH-1:0] out_7834;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.125)
        ) inst_7834 (
            .outp(out_7834)
        );
        

        logic [WIDTH-1:0] out_7835;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7835 (
            .a(out_7834),
            .b(out_3),
            .outp(out_7835)
        );        
        

        logic [WIDTH-1:0] out_7836;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7836 (
            .in(out_7835),
            .outp(out_7836)
        );
        

        logic [WIDTH-1:0] out_7837;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7837 (
            .a(out_7833),
            .b(out_7836),
            .outp(out_7837)
        );        
        

        logic [WIDTH-1:0] out_7838;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7838 (
            .a(out_7832),
            .b(out_7837),
            .outp(out_7838)
        );        
        

        logic [WIDTH-1:0] out_7839;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(3.475)
        ) inst_7839 (
            .outp(out_7839)
        );
        

        logic [WIDTH-1:0] out_7840;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7840 (
            .a(out_7839),
            .b(out_3),
            .outp(out_7840)
        );        
        

        logic [WIDTH-1:0] out_7841;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7841 (
            .a(out_6858),
            .b(out_7840),
            .outp(out_7841)
        );        
        

        logic [WIDTH-1:0] out_7842;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7842 (
            .a(out_7841),
            .b(out_7645),
            .outp(out_7842)
        );        
        

        logic [WIDTH-1:0] out_7843;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7843 (
            .a(out_7838),
            .b(out_7842),
            .outp(out_7843)
        );        
        

        logic [WIDTH-1:0] out_7844;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7844 (
            .a(out_4175),
            .b(out_6462),
            .outp(out_7844)
        );        
        

        logic [WIDTH-1:0] out_7845;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7845 (
            .a(out_7844),
            .b(out_6477),
            .outp(out_7845)
        );        
        

        logic [WIDTH-1:0] out_7846;
        const_element #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS),
            .VALUE(6.3)
        ) inst_7846 (
            .outp(out_7846)
        );
        

        logic [WIDTH-1:0] out_7847;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7847 (
            .a(out_7846),
            .b(out_3),
            .outp(out_7847)
        );        
        

        logic [WIDTH-1:0] out_7848;
        fixed_point_neg #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7848 (
            .in(out_7847),
            .outp(out_7848)
        );
        

        logic [WIDTH-1:0] out_7849;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7849 (
            .a(out_7845),
            .b(out_7848),
            .outp(out_7849)
        );        
        

        logic [WIDTH-1:0] out_7850;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7850 (
            .in(out_7743),
            .outp(out_7850)
        );
        

        logic [WIDTH-1:0] out_7851;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7851 (
            .a(out_6498),
            .b(out_7850),
            .outp(out_7851)
        );        
        

        logic [WIDTH-1:0] out_7852;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7852 (
            .in(out_7851),
            .outp(out_7852)
        );
        

        logic [WIDTH-1:0] out_7853;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7853 (
            .a(out_9),
            .b(out_7852),
            .outp(out_7853)
        );        
        

        logic [WIDTH-1:0] out_7854;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7854 (
            .a(out_7852),
            .b(out_21),
            .outp(out_7854)
        );        
        

        logic [WIDTH-1:0] out_7855;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7855 (
            .a(out_7853),
            .b(out_7854),
            .outp(out_7855)
        );        
        

        logic [WIDTH-1:0] out_7856;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7856 (
            .a(out_14),
            .b(out_3047),
            .outp(out_7856)
        );        
        

        logic [WIDTH-1:0] out_7857;
        fixed_point_square #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7857 (
            .in(out_7856),
            .outp(out_7857)
        );
        

        logic [WIDTH-1:0] out_7858;
        fixed_point_add #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7858 (
            .a(out_7850),
            .b(out_7857),
            .outp(out_7858)
        );        
        

        logic [WIDTH-1:0] out_7859;
        fixed_point_sqrt #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7859 (
            .in(out_7858),
            .outp(out_7859)
        );
        

        logic [WIDTH-1:0] out_7860;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7860 (
            .a(out_9),
            .b(out_7859),
            .outp(out_7860)
        );        
        

        logic [WIDTH-1:0] out_7861;
        fixed_point_sub #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7861 (
            .a(out_7859),
            .b(out_21),
            .outp(out_7861)
        );        
        

        logic [WIDTH-1:0] out_7862;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7862 (
            .a(out_7860),
            .b(out_7861),
            .outp(out_7862)
        );        
        

        logic [WIDTH-1:0] out_7863;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7863 (
            .a(out_7855),
            .b(out_7862),
            .outp(out_7863)
        );        
        

        logic [WIDTH-1:0] out_7864;
        fixed_point_max #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7864 (
            .a(out_7849),
            .b(out_7863),
            .outp(out_7864)
        );        
        

        logic [WIDTH-1:0] out_7865;
        fixed_point_min #(
            .WIDTH(WIDTH),
            .FRAC_BITS(FRAC_BITS)
        ) inst_7865 (
            .a(out_7843),
            .b(out_7864),
            .outp(out_7865)
        );        
        

    assign out = out_7865;
    
endmodule
